��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n~����1cg�&Ft��ͽثc��N�i\r���y���AKK^�z��U��Z:�;��KP�B ��N��A�>	��h��H~,
�z�*�M(�b	������LV�laD=tp8F�+����Rq�����������+�nS�U�F7&���S����"�M ��U���@�˴�5��.� -;P�~�oa|
)k���BЖ�@�o�v�4ߘ<��4�l��D�4Ak���-.b���mC*��D�i�M%��%�k�~&ʳ��0!����nY�qe��3��ck����o��z"��,f�ը��%$���|�;+#�0f�UhOǃ��2刑�Lc�����|��|����Q��Ol�pf��\�4Y�
A�Y�a@��qnNAz�pד��ݮiF�?��'~&{�X�v����H�	���Gʲ���dӤ�>v�� ���K�B�x��X�[#s��W�V��.��f$�n���:Qn��24"M��<48�}[�� �(�5��t�L�6����ئe3Xa�|=�X$nD�H"ď�Vl��⼞=��5��n�Q���6;#٬"I�L���P����/P=�}�㟂���C���?�ZI�r�	5��]%���ē�2FTC�Sh��Ds]鉬�@�0:�?"ܮAۙ�>���?��i+c��$�vf�:��P����LX�Z��+�'��Y�}�G��)��q��ʋ�X�]���ۅЅ�aڴG��i����(ް?	�P9���y�
�����E==6�iS��=م�gU����!��8�د�§���g��d���B�Rx%��E}��8�!-�U��@=�R ��s�/�ǥ�;,'�f��|�<�\W�21u�a���{-��������k�����@b��G�9SK{[O��Y��7�vb���yS�����	�63ǲ�Sr�,B�/�t�(��� bc";W���"-�����?�1\�ؤ'

`�x��4Q.�H����E�l���5��S���kd1��{+Hڔ�խ8�|$�������؄+����)���gn��+砯y���>3T��Xw5ӗ<,�C���   ̰�78ys
7�s�m�MO���_���t�3���d���*�۱�)!܃�9��-�J���.��qkT�*)�
0�Fx����t�g#@p��s���(��ܐ�q��U)ײ�Zƚś�!����qp� }�̚�5�*��%�̲[�����]�c�Sk�}vvIw��9TY�WXWmd͸��ל�� $�	���Ʀ�˜͖�"���A��P'�k���"XT��O�荺���UÁ�jô!���N�΁F�\?����&�5/��B�xAW����'��GZ��P�qnǔ2Z�����ے�@�/͈���S�Q�s���������)8 ���RKW;�<g>�X|��E�,D�~�^L:A�[�ߋ�R[\��=�IHDѝ{��=A�Y���X0�N	�_�x������?���ů��q�շ�t�0��R��>���m��'�����c�g�?�X#����.���g��B4�c�/�H&��^�l�nUS,�N�"N;����L7z��/A�W�ͺ���&�pQ�q�`#��b�c�O_~OP�	�����AƝ��.�TN���-�Oc�������c������lP�*��u�r�J����3\�g"���LUH��6%��gJmw��y�v���,(Ǿ>�*~r�[eX�1���}G�z��c��?�{\v�����W��e��Wx�h�>$Q����`
,�EY'�<9`���17Z"����a�3JMb���*-iͶ��!Rt	6Nf������ũ��:Z1�����i�-~��:��9Ӊ�N��LL�b�$�Ę�/�� �!�̜}in:��$�g0h�\�f/[$�$��B���-g
S��o��x ��a>WEQ�ZԿ�0��r��|[���,�ˁP���p��b�^SP�uo����}3��}�;;���l����RE��h6c��/6��⮍���q��5)Q��6h�Ѳ��&�0�Ą"�늊(��^�n�)�����gs��i({Su�&�ռ\���H#�ǎ4��X)]�c�ꩻ�R�Q�
�Y�a�U6���r��V�����r�	��W�����Ԁ~���?��IH�\0���y�ΑN�b挮9/qT�s=�l��~�v-�r��oK,Ă�Z�I���W�G/��%���'�U~ҿ0��D��r(S�eJ{�5Aw~�蝹!h	vu[��Q�?-2���n�Vjh�@���ܶq����ywT	>�߶��/זh||SHqb�`ӡ��fg��C�0$ o��w_���c�x���7a��1��Uÿ�*�Q0t�����~Ȇ���5̤��Μ�nbP���{���@�B�5l8���&AR��󮻴47���6Ӟl�ӑ9��a�[P/����XoHv�.`�3�*�x�6F�yI݉�C���D�*���-9�'V���%�ޥ��\M\t{ji0�Q�Sn[���j��%��~~"n�����bI�]
����p�gEYM��Գ)�/���=���g�z:��ݷ$� %t�ל
��%J^��ЎUn�-��1oщ�,���Mϵ�+����S���ׄ��'��Y䕷���l�`���z���5�,�]��l���Y���H8D�37��ϐ��O�p��]�N�-2����J+��X��n��aaU��>�����P���jaX����3V׌M�N��P�9YN!�q�yȶr�O	�,�/6�V�$	�;�"� ���1�s�]��4�к�{�M<�^D�o>=-&�[����b�#(p���=v�#�8d���p��C
�� (_�Պk7��Q��
���s��K��K<UF�5�P�Y��.|�PC���l�E�(�Ojr_�R����Q4C�1�2�g� _�P�?�5�k����4T�iS"�%̃��g���N � I��8������M�Y��#���|d�~�ҔMlkrISc��Ÿq�q;�V��0���9m�!����#VZ~����︖��U{x`���܉p?a8�}O�3��d�.�^�nbh
�u���u�-�a�:�\@���!˒D�9��sH+�I�x�������?����Y�Eq	�,����f��э.2l8�E��&[����J�*�ߑ�-Rq�,�G�//�2!s��Qik3�)���T��lH�tYT�.�HV;*��$�{��":�\-P��~��+�ì_�F�F��:v�T�S�Z��w��"T��Ĝ'��C8{�_��h �)�6n���[���Ci�~�W�O�Ԋ|�Q�T���&� їnz�XA ����m�M�*��+�q���}��6�خqSR{	co��~8~/v*#K�^����������U	�G9��Wy%'��M���a�l�U�k��� �y���=����ҧ*�^�k���B5u��S#;�d-%3�sY����F��>EC
WCC�x �P�ZB Ԉ�!�`|Wc�����WC�w��ØZ���NX]��y�-7Q����^�+���ʑq��Ѭm�b�B�O�k1u� ��l�0c�I�����č]��^��U}Pq$z�b�ɭ"r���C=��Z_EBD���sm.�E��=s���iA<l'�`�e".��k^�z�<�[������S���K2g��S�j���ꔂ�R��bH�0���8�<�S�T7�G��6<Hy%��Ȗ���%��~M3��p�%b.ecM@����/ezCM6[+�-�䢤���t�LI�Vh_�hrNS1�R�^��ܚ((4I0ڃ�j_��K�7Iv�ʕ���06:wIZ�6�����Lɺ[o|��}���\	&��M���I�[�8Ԅ_q����w�\A��y��l��-���s	����6����:_���w���l]b�gM�ϼ/����O.��r9/C�s�`�Ő߇I��"�gW�ג +Wⓘ}\���nw��%�?�a�D�$rJX�_on��Q���"�j��q�/��a2(`�>�Y��k�x�A0_���0���D�HhiT�S�5dǾ��yǽ��3PP���jT����n����9Y�ѡ>�(��Rgfs/�������f�[lC8�$%/B ��=�-E�Z��դ\�>r!2W����1��&8���� �.�0�H�m��2j�����u��#3g�����Z�QϰC���+4���e�9eF�͂���z��zx�cb��z(�ȫ�Z���
��%�V�#t_1[8y������Մ���QS�{7�_�.^�LR�����=�_<��U=ψ��%eο|?���]�d��E0�=w���jR"����ط?vN��W'�l�	;b��L)�<B��&BPy�t�Wy�؂#�k�3�[�-��0��h(�>��ӿ^�DA'׆��a���ԧBM���Ao�3��w���@,����k�<c8�,�yF��s��}��Kz�`�0ˀ��h�V��0�^?��S0:��<�Л��A�X���1�
�$�m�i�>�V�ۘ�td'��Kj������U�k��g-a��K)�Q\+�H�E�zp� };(@Q�����bM�����LN�C�:9�6s��RO��'��"AG��󞎷碊��_��cV�V��I]�fUE���SʚR�Ǧ��i�F +݈<=�́̕:�Ѥ�^D��'x��x���^�N�6���'b]��;�H�Q��>E*�t��%�:�1�mD�r���ex,m�c�@x!0~�q;��r��"����5�ᠧzz�l`�Y#c݌G���kFJ-���Q�V�f���z�*-��&��<lD(v�;+犹R�����S�6�&bM��������t�G�	���]�D��������pZ$mYP�e��.xM[]bO��|�ϱ����k�_�S�_���e�[l1���T=M�
��?2��t%c	Z�3[���+�(�,t>Q}��9+%�`�q���-�J��am,H� u�+�b����W�-%nҶ�o��/�V=�H��7ʚ��ERFI�|%��mNBX�6~C\i��]�: �l;	�ؓ��iSR���oT�z%�5m�I�jjxqݒ���S�
0�ϱgҎ*�G`+�e����܂6��)�c2nW�b�3\�M��v���F��E��y}}�x�!e�Þ��p!g�⁖�A��D{oZ�	�n�:x�o�d��Q'�a�Ɣ��C4�b&E"5���M4H��z�3 ��W��ބ�W�2c��26��4�^�tn.��dώ�e���Ɂh�EL�e+����d[<[�Dv!��Hh�?�O�6�͢��Aރ3{�Op�ҽ��`���\C�R�O�1{��W�����r]�7�98
}� 3�N��i�>v��R~�*�fj��da�vj[�.g�2�&�J{��`h�I\.��h-=[R j~���ژ2�Q*d��nΔ�uEv�����	���7���ae�s��ܻ� �UiX#dJ��y'��J5�u�4<�(�b�L����/)?�WD�د��*����	AiH@yiJ��5��)�i�'�M�~9L���_˶��
�~!���b��z@dD�{�n�r���Q���|�t�;�!�P�m�΋\�~�ǯ���N��Ⱦ���{�:ֳ���/F��r�
���������(T�G�ύxEb���/���øf��Јdtt9�"7h*��#;.�Ԣ���dS�1�@9_bȸ���d��y��a\�u�+w�* C��W|a�S=���"��f�V��|@����rA��`7y�-�*���-J��.X��N�TcL/�SE�A��e:B`̖㬙��s�{D'�p��.�12�$服���g���'�^�()R^��͜���γHxH���w���4��ņ�_z+Nc��I���2�EL!P=T�x�˅�\Ԛ���=6�Z�բm�S�:��"u.��,"s��s�my���r�b(W�H���)��	A�"�Z�΢�.�L���*��r3TR�%ww�7��2p�Z���%�����L�Ro���<L̑�ZԂ
�� G�ۇ�uc�i؀i�Uۈ�ݪ�@�ǅ5ԣIJ+/��>���ICh:�5L8&��I\_�1�ï��˜A)[�	1=��MX��Xg����.��˥|��VQ��N��0jg|���}�]D$�Ø������D���*JW�*��g;[��-�6��S��Ht62d5�e j�\u�{�9 ��	PBU�e��/<��dIU�}5Lc�_-}���E���g�T��0�.�A`����f��w	�����;r��r=kb��wt(ԤO��t/��X7.�'rd�Hh:i6���yҺ�e)awhKA�.�N�w)���1�{��f�b��7?-(��=s�Z"
B�JfUdR
�̔G���;�~�W"�_«�Jq�}S鶩����z$��jM�����h�;\+�����cZ
�62�������??�@��X�W�d�i��m���}Y��)�����n��.xC�ŏ��IRt[��Π,O���5��-H7)֋�����c�#~w��2g)]f0�*mAn�@�u�v��#5��g^�,U�d#��!Bd����_�wz68�P?��^b��n�A�#.�0h8��N�\�`CBR�Z��M�26���P�t�R}�I��+�Z;�t	�Rb�?�~CB���nd�־_k"�H����&�>��q�;�?	k�H	����q}:�)ȒM�9��}���:��Z���������Qv�*=t��,�e8���Q`*@��
��Q]�䬑t@5�w)�#=om��j��R&�@�&�oc�@�Um�6��RX��aw�f
�bm��O�I�U�6���Ӵ�j�LI�wL0�N�͛ѡÍWurY��/C��� t	$���Z�σ�s���S�Tb�Dо�����E5�}}u���d��?ۓ{����p�k��M��9��E1�'���q#{�|�Q{��E��ᓑ�4;B��/YY-x1��Y���Hx 6 U�c).{�|��5;[�䯙7΅��ٱ;Sjz9�G*�E���h�4�/9%�7��g��~KK���W�e�1�m:�\~3*Ov���?�qZD"�a�>7�r(�N>��>���O�E�����2�֏�>q����6e�7�T��M���=ȹ׋�+ݘd�7���#������)R�Ĩ�6b��md�e�Y�n� ��3eM=��'��8�ȉZ�	O���`�L�d�n���*c)jp�^�vqB+��W�(O;aoM�ٞ�y��p���"˕|;`���PTl�ǉWY��c�%��n~��0��j;����)����N�&ԖwR��&j�9&��Q�+#jHxC/�e���p����d󨠘��NՈ��*EV�9�سz�L����kV�����] K[�)+���.����G֜?\��_s^g�L��Nn&������'=}��֒�kv_�uN
Ф��+��\��D9R*�=��rʂYp��)Y-�Wm��$���&g.�ʣ؃y�����h ?�+��0��?G~i"�$���,�kY, �y�)�1 I���v0Q�t���^��q��W�ajV�f�ڢl&�k���U7���;a��m=y� Q�<mo�4r�6�T�,�,� �+��1���6��'}X+�h^�z1����X������֩��5y���46"���Y:"1��,�����k���*-g��lV�g@uލ7���Hbvb(�#}c�w_�^�"�(���e>� ��X�������[*�pɹ=��ؙ��5ڞֿ�Yi*�TQ~��؈�茞Dh~4��P;_~21�݄���l�I�O��%�t��-�%Iy�ut#�L�<���˽{�`�	�6�;pږh�3��:�O<WsڻK�Dv:�t^uѵ���m��͐!BN��D�)(������>u���bc�G1G�Ň�j��,[����퉻t�f- �y�:��܌��!3��` j�Uo)7�d��ٱX�������F�]�n�q��v/L�_9����� ˸.�h1��	�T+%����v|�\<{Զs�O��Le"?�O�Кs�1X|Q��ݚ��.h�:h,�ԟU"���ȡ��\�v�`�TW�}�a��f�9�KS�>��'ڒ�I<&h`�%�I�)�Í��Gm/S��N�[�2�4[3(����u�R�7R[�3�&[Mvl,0�Go��#̭tG��yu��HК���36�q1QI�d#KX�p~��o�}���䆗=��I%<��S�\c�*��V+��%t;��|�H�U���A������)��� �[������A{�Q�&f ���(�i�y�{����O��%�P��}��憕2�u���)^�si�Iw��ԡ��B�/���?r��={��ʀH���)!X�P��A�4y>-�K��r��s���X-��c�|���D90�u���Lo���Xa��{�Đ=��� ��1*���a����~Я!h9�"��AyB-b4b+��m��Ol��d�=ɣN�]�W�y�1��P15;�=���?��y�P\�������ȕ��ØAQ���ߪ���}R�H�J���'8����-�ԁ�t��L�L�C�G}k���9�xi�tM��a�k�dl��C��Br��_��g}�֠7�g���KJ����{�w��t7D���/���]�V��p�H��xq�Ж�58W<T�ٌ��us�u;r!߃"�'����b�$�U
���ʗ�����r�̛��n���J4	�UV���������!̓XK[#o�r'
~�Y��ut!�F�[G�T��ھ?M�t�Jӟn�f��l)�k`��U$����֯O�s�+�r6�a��'��~ա�����["n%����f��쉦�����t3�D��vG�7.�iE�a�����!߫ZV��1����Dl�e^�,V
����x���]D\���g�f��`��n��J�]{�f��$w*QY.�@�m3~�Z�kW9��Pѿm-���L�?�[r��(Fl�.��{�$��9��Iי�?>v��K.@B���hAUQ��X�8����K.He+L0��H�;�9����RZ2U����;�,\(�	
�g�AG� �j>�c���犣� �>٤񸀫�xu�.AJ$���cP���?�i[�u����D]��!�U{t�Z�u��X��ǚ_��>d��뗆X���lo�y��IZk��ٿP,�>�e�!+�m9�EV�Ǔ�e�h����{���������`e�ۀs{���#MC�z���g4ldU��@!���鸙�*�%�����'�:�~��r�.g�$u�d��cBԦ���f�*w��'��4�$H��Q�׽<˲J�����[�Sb��7,����o>*��=�y	��Y?L|���4e/gQ3���� � ���{�f#Ҹ�M����5[Z�����D����Y�i��R����#5#,��弈�IE��X��Ttύw�R��\�Yn�V���	R~�����XwP � w \����ߌ�p�Q�kb7t�k'��$0�aL�g�d��0�cX��Z��+{e��囂�mz='y�M����k�1/T;}��~s�)s���wh���	M@�U�)6��N��/E��E}�rUX˫\q������phP�I���>2~�f_��EEs8rl�Ȥ87e)�RU��ki����;��Z&}L�.�>�[���,�I�z:�}^�X�DCjj�\�ȥj�f1SG�P�V=�+f���b5�&$����Q�����l�����*X�u՞�T4��%����p�3�fqy'\��f�p^�*��:��Cl��5X_��;|YL�tG=�}*A�]R�ټY��҈gW��;��a�7lm��=�H/���L�Z�g ՘f�C�,e��~�/:�'��X����(��(�V$7G�)��D��oT���jɥ3C�z�f��|�.�����6X<hjC�F��%%�!���>�g�Q{�({]���X�A[>���z/�u�q� |�Xs���ٟĺ��_`@���`C�}�3������C!�B��ht��bn�}Uʡ��Go�j��#sbES4W��ǚ��Y�~_q��J]@E{'�gl�)����0ƶ�	� 0BL(�+��f�5:3Q�t�ȸ驦���Lb�,~���"���e�SE_���x!��=�bH���E���j.'<�W�w��]�q8W�Z��N��a��⫒Hd��5�7�����g�Zy��o�F��W�r��,Gᬌ>�ҊC�R��
��#E��+`�*��V���u'Q�����U����&��=�?q���l�7���Mcv���Q���m�����S�c��;u���Jܢ��5��r�cO+�;Q�V�Z�����{*�1���Q�Wo�R ��)b޺��e"o��^\���}W��'�8�;��	p�4�,-�����X�_�En�R �>#N�u?�XIE�ٰ�q6��*P���=i��^��e�YA�C7R.{��������M�݈5Pw��T�M��tY2?�>`@��B85Q����.
 |ԏ��Ez�I~�B�I��#����W��6�cd��J�w�6�'�!�ܶ���"��"��{��r`�U�rS�}o�h4%>�;uc��1Hd��}��(�
0�p�6t�}]������p��(�Ik}M,G5���|%m��jg��(<���;x�_�`�x"��#-��|a�ƹH���\���C�h�?�;�fLd�"��V,R�-B�W6�^��] ���,��%�p��ZN����=�1<8*H;����P��=y�2���,�l���R�y� yo<)j:kC�@���wN��"��T0	��~U�iN �p���k�5��8��"��GKW��XKF��o�QKC
[������/	U��Ŗ��g��W��c���I�'������6�K�l����v�u��������8"n��AS.���o���5D��i��p�YeP	}�2�A�D)��������y��(	G�ܖ�0%z���Q �`�� Ϡ�
t/�U��Ҧ��#sX<P��Z��i�\�p��|����o���2����M ���ç��M�z1(����Ә�n�Ub����h�M�}a#���MyU5��F�s��b�;x�Bį�A@Ύ��F8���䑂!w���D�VP(�4�Y
����k�5��ԅ�1=~�i�� �w"���*���CZ�q̈́��M+s}��M�)��U���3��3�s�ӿI��P����k�W�c���ʠ�jn�.g�T�=��ƪu����>kʩ�n1��Ӳ��6]��(~r\�p���M���xD����Ũ�p|-/��p��ԧ��=�tA�2У��Dz}j{N�U�(�*����Wsr��9R0����ϑrd��Ϭ���^KK�$�e�9�9�Pc!�^���+�.Y�ߑS�)�x{{d^s�k)}�[����u/L-�<��0���MQ��i�qY�L��@��<�Z�+y/���e>o���D�M����(R�ETX>v���`մecV$9�<��⑎������+V!�YYz�JH7R�r���QEǈ�w����,�N;�������)����P]�]a7��yo�m�}*�	�Y���%$,Dz�'� R͕,�;�N1��]��*���k��zϦ�ҡ߂�+�>�vfܾ�J<��%��C&�P`~�/W�1mv/F����cE\+X��)�v*���'�T�Ǎ8����Ѣ)P'��L���qC	�,�poͱ�N>�~��X�z��\eo�W�"f�Ժ����_�K�nAm�k�#�ȁ���ե�}um�(&�����nO��Kf�|��<�+��)�; ��	8D�򚨃0Izƅ`���}�v�pmm�{�F=�Z�@,��P�ъ�d�IB�g*��Q|�s�u^%�G��E6��ujn󺎜J��=�r����aC{�	σc��-])9��(a�H��1b�6b��e���\R���>z�aּ��?��Q"��� �ט��vƕ��t�f!*%���5v�T�����*���|�7v���Y)���N�(u��	ȿ���&xLy�\����D�'��b���<T����Hv)fo�MJ�n����*��DO��{}c ew����fϤ�?�s����E�(Qd�hs�	w�X%Mk{ض��at�5�Ҋ	�̌L��ڐ�����P^O��\��} 40� 4Z�e|�A��/:T�.o-��9
�7���K�B��:��<��������o�X��=0W��S,z(�_}_��C����3wϭqӆ�T���lvҶ�6$}#~��jͦ�H��z��P<�v���;����*w;İ�����f�+;C�����h%_�����ʈ�*`��S�?��I膏��k�����$�
��h�e�_�g7��i�/�p���l�����>
�a��d�+Syx6�u�4Sg�D�&��Ҋm�L����O/G����g�Aa<p��#�<�݉�p=�Kn���
y�	k��(J6k��mV�-n,H"��J�(�!-�^�J�xW��x��B)��'�]@{�1����C|�N����?��h��*��3�LM��Aߥ��R����G�8��R�2�] �V�4S����W�����N=m%�EM��4�]W�0:fR���C����*H��)�̂UA�]�T	�P�7�[��<u'g�`�6���4���Am"��A.ib�{Nw��vP�����
�������_eb.�^X`53�Y��ह��f�a�����v�ʽZ2���4�mK���&G�1j�k?��7���*ZL�x�0><�d�(s�_��d̯���c��(M�6�5p94G���}z_n{��F��K,u"��X�&׆���1$���4����E{F�!C�2��Zy<����a<2�Ӈk��J����b��ib����	���U\��hU'L�u0۴)"�:Z=��,�m΀V?^�ݰ����{7�9�)���o�G�^�,,�#����+��jE�I闂���SJ��D�I�h̪�k(�B��7R:m�a&砧�'lq�wC#~@'������m^m��K�"�t9�b����m'�Ї��P�Ad:������9G'�����Be������j���b�w+����G�p׬f-�F���3w�A���S9���l�n=.P�&�}�*g���g/�Ӭ�2����n'iJ�}i3��N��ƅ�Y������b-a�E����Xu�A����*P���c�aZQΖV�i2I� ,����}����vֳ�:RN����h�ܥ)��!0�E�7�6��iN�!\������5�R���k6�9�Q��1X
"%G���D��6��eM���h�8�����ɩB�?a�U�ҙr�=���7�v��T�}�X�����T7�]�����g�X��ӿp���h�Fq&�iJpM�r�.a���^A%��?!=��D���a��ZmR���d�r�T��)�d^�Ԡ���;E�a&�uC�%��7H�'G�3J��r��do�N+TӐ���;qvX�ڦx�)X	�_�;�J.t滠���A)�y�N�<�����W�va��⮰p�J}YI?�X�~�V���Y*� �\�|/B��%qf~�mR5}�S�0O��?�$���*薕�Z�<\J��`_]����z��a��D��2�wݯ٨�2s�Z�m��-S�z�l�wPY�4��-��zN�������f����oȕ ��R�	B�=Ӓ����������>��*�.u|�p�ɶ��N�n&�/�do1���xP����s�ճ:����νѠ����z:�o�ćnF�+k�{�:ڢl�A������H/��J���|T[ȖU8m%������@Ѷ�ƹh��-��k����ϯY��a5{p*`l��Q�?�O��z��0��^v血�cfm��XR�1�2�  P����R�N��|�qCaE>Yj�b��
&~����o�ۦ�9���s�1���X��d] S.��Ǒ�$p�R���RW�;��׼S��~�q-)xp{�z���E+�vKM���C���n��5!�E��dx�(R�U0�P�PE�S����|stA�^�"������m��EJ)������"C�[�F���+1�����yG5Y�o䧥�8�?�����p\G֦iUc��@琈�A>vH%П�G�@j���^0��9C6�[e��;�_϶ד��0o{����55��K1���zi{3����I����Sz4o�>y8���R�)v��*��R�,��^;�;�?�r����w���j�h�R�ֿ�۬�/�#P����P_�c�����·!ɭ�j텮E��W�s/" 㡘�ފƖ�|�mʖ�9����H���AU��Χ�1(q�4�r��4�P������~�9����U�������{�e��rc����S���� ������뙫�p�����>�H��d�7�RF��=�G�:p��/f�/�o��D⏥J�q�N6ȳ����"��޴u�sa8�p�Wũ[�*�_�9]��Z!#�L���yw�j�� f�Pho9�[�D�D�6w��IƱ�i����6f:�L�����A�yv�� ��A���&�ݣ���@�-8V�$��$�#-j��i]��;6EI�&�]:a������Xt�69n��P *�̛t��xAx���{'L�v�|�Wd��ϔ�&��w�uVOb)pu�pL�U�џ
Ϟ����~\J�^�s��Ͱ���[P�(�n�&��w�Ҵ�Q�3�G�-��X�Q����R��>C=�
F��	����t��Z E��m?��^��4?��� �0R���(����;i_��M�	4��&���R�����������&raS���)*����.i��Z�>:SUy�Y�H����f���x�;J�Xg��;��b��b2�N2�4�U,סyv''^�(�xh)p��pX4���Y�߷����y�oL��iTͬ�����L�ĵ�0��,�:��������ڣAnC��Ѣ�.V�)��j���e.DN�"|�>ˤE�����|{�4�塠�:;���wg�׆{vp�k��`䆴שvqŕ�eG@a�9;�%�y����y�1:�����ہAO�p�ǘ����<��z<�h�c�r1����AgW�P�n���jå}-�\bм����f!TT�����mD~]y��f��	�W���h=:Z�
���4�ݖݓ���*� +wн	�t��>��'4b���/y�ɭJ`�	P/�Z�5�m%�	уcIV�K��,g�N�5c؆�f&R%�����R1�-�Z
Rd/�&OH1"�m������R���^3���9`-N����2N����I�N�	�l�ŃLn�h�1�+8*xK$4t�̢���(��b�MA⪍��\�41�y�T�M��D����w�����6��b�Qo2�xqP�	�s��������d\�# �GH�vɹ��}^�Tt�*�-�b�����֬��&k�x��qΜ,��(�<c����	]�ıˣ>�Y��_�2�UI�S��ʒ�D�%�S+�*�m�\cS".�gx9�R:���fz�ü�N��(K�L��H&�A���6	g��n�CN��-����S`��x�ah�W�!r�̓��]{�w�1��r�jV�s�}_�:�3T�W���Z�=���(8ڻ01T��꠼߮�	�ʴć���@�C:�&�b��O�J��K�ZB�R���ݨ�5�j�輓e ��G	6ZFtw����ߒ�l��x؞�¾a�y��>���apmZZ�&f�h��Rg}��J~�������g�;�:�|&8���ƫV���&;�6tC$"�}�X�KL��'��̧5Gw��qb�V�����K�ƃ�R���p 9�Z�$Y\��Yv	�E�%�����*G)<�&��$,�/9c�$����wٞH� 6��?��|�AW��͓=���U�����Ϻ�b�Rm�۝JX�Ș��&�SC1�?��N{w|���	�&w�/��N*��'���I�ݷ���/C޳�F�/?)F�8�����%@�1���_y#�����	��G��}�\�W�7�����՟�4Xc�8�;��%��F����v;�j��j;N����5�D�����������:�tvmjͩ��',/�`���D�U,���I��/���ƌ@�c��L��6�bŰ����Hג= ��!�!�o�����B�N�5��^�D��0C�7�+-��ҿq��'E^yHO�d(�j���k�&b�2ddL�]��(�{�2|��kH`��G� /��VU��l�z������T�-?C<;[�Q�iFr2P	���=Ɋ���������EF��B%8��t�$���C�3� ��7�W��l�@v8���1�x�L�ǥ�֖m$�2�~�re5�l4T�|����$�ϖ�5䍨��{1 N�t�m;ܡ0A�Հ�	�	p?v�o.jn%����� d����ʄSJ�І�Oɐ�n$�gp.R�h�����m��|t��(i�p�.�PoO��w6��M�=U�0X��6�@%��D#�:dV�Vgq�"�9$���ؑg�XQ�Tz���9[���hIs��-�|]�T)���k8Ah��T)X��Z����D�DE �����gǺU_U�F̏ab���Ƶj�B��#F����X41��Z���z6	@.~
M��e��и�ܜ1
++�h��V�g��S�g�õI����u%�2����T��c�X�8uݎo���W�&�C�}�fl\2�z�j���������ȇ:~�����
i�]�jL�������1�
�5�<�%��7X�r�y�%�:��B
x��Qg7����m�[9�g�!������C���c�]�+�0�ɘy^*!��$5���K%��aw|`���k-�wՈ�ϲ u?��r�c�55��j�����
R1f�<��~M=�D��Vc*��B��/�4��J��i �]3��e��pM���R��n�ҟ6�ʺ7�$���yR:�`��d$Σ����Y��F$}@xv�a#M,s����X{"�s��&��H�s����3����H�%����/,�}�iV���v��z�|?�}`P#"�MeDY[�Yaկ���;�I��c�f�w�?�!���ER?Xغ��X;�OC���:Z�Vl��x�]~ŌڇȆ�p��A���p3~�GF�ڻ�����.�(��0Ml3�2�|��*]���e��p�~r�l��TD�x�q��ftu�E�hZw�(c�d;����Ѕ_���l2	�k��_^1�x���dC�sOQl&�VvQ� ��w����e��)�2��!�m��u˵����_kT�O`H���$�ū�h.Fk��J@��(D���W�Lq�Oe�=2��b)�[�9j�a�}ƿ�"����U�k|�,��� �'���4�\� >ԨHz'aE�^ˬ:���w|�)>:���^���!����&�x-Cb'��p�l�ꛘ�fͥ�F�V�=�P�4�)꽗�A����ï�b>c�9������W���DZ��Eڵ'�o�y� e��-�3w�Px��H��H/u�`'�^gJ�2�j��h��>XƔfljJf�Df;���sn�o}�u���e������c	$��DgYɄ�vA�C�����;���T�'[�ş�C��7�AvF���#3�,|��x�+�ۖe�'ਃ9nM�Q�Ѥ�1z5s�_�
Ԥ���0��u
��,\U~W� f]v�ij�c��tj�1�=J��w��t�.�Yr;T����.I�����F�v�_Xgx�����2vuܖ�|EMAi uw����'�z ws���,���=����S����j��L�C��R�ce_p@��<i��}� ��u�P������H5��+I�~s�!� �b�Ǒ�E�w�Ә�0�8�2��#�P� Qz�T0=ase�<_�O�%�n�����ׁqo��VhRr2�K~��o�����*�)2	�X�.L7H�{�X��~�MM�5�������{�3!�,p��|�����?a3���z��9^g���iz z�~$�o�>�wJ���I����¿�,��<��[��^���17@;�B�1������[�ʖ�	����G�
���97}ޟ�t]��#V�/� �]�701TYHI�H��B��᝘��к��2;�伉�qq�m�J�CYа1���DB:
BO��;J���A�FAu�(��.Ln"�ui(�Ş�>�~��<���e�N@�-c��V� %c��N_,:]r^k9p��\,(HG	%��hjk�V�8��p��gGG� "S̋�N9�ϻ	c�O�q�.�L`g���9P��Ă�Mf}���
C\��hS*`Z���utK�a_��z�1�Ze���� �u�3��w�]ĸ�F�	ߋ=��.��+:@�`pT��J��2^�JS�#����A����;Y�������Nk������#�!���ԏ��(��F�;�PG~���=��<o��[��~nP�T}�*W�����j���![�Y�̒߾��� �R 듹�t5�]�j,�81R?��.�Do�vj�T�un�� ��w��:�_�v*J h;}�.D�c�8���G輫���Jt��.0�vqn̒M��^:�d���ʪ��y<�j���7�Ǉx�_������av���w����?&�=���I�Ǩ�0�q6E4�̚�"�U%0���GR�~J�Nϲb��p�o[��7����		p/���	����t�^?������$�[�� R=iɢ�� �����훋g�Q�\y�3�p���t�( p���A��}-^c�J����b<�9<��.6. ]�0���`s{\�h���+k�b�.k_J$\�Dl���R,��g�!0,J+�`6[������XV!>_���K�.�Jjg�N���W�(Á��qZ�q�vP*���'d��ݞ=]GPxw�7xR�-&�S�z���?؜/���N&|���[$�;u$K�~Jeg�0�ՌI��
dО���7��(m���m�\`�}�樗���/��wiI� Q��Z2�N�q�O��u2ytT��㨈���W܄�<�IN�߃�݈q�F�̬�ɘ�1�iժ(iά��;Y�����c7�H4������'�p	r*v\XF�Y�< mT�A'���fmL쏡�Yb�?�JP��[9��u͆Cd�cO�yH��W�׬^�u���C�+�:���9�$*�������lE�r��f�M_י`��(_�+!)�!�j�FTr���;�q��$�ؤ\D�J���q=���X�(��H2�b]_��0��M�c�L`R�҉-,�RK;F�����j�0��n���a�;6b�Bi+1��������z��Ug���d�ދ���O�_�=zx��m��7�x�%�`�9K�|>
mPZ���'J��D^�Fo�g�IV.,�p�}�k>�C��])�7S+d�W�S�� �PcB.�q�3�ת��K������^�m�[�$��[h��=��ijI>R暻�0�-�L�D����7��hk���W�/�sj��Ѡ���-��̃�_��T�^���C�q�J��m��ؘ��N�pv.�+��~�FBV6X����s���T��,47s]Ǝ�@g}t�%�X�v�ҩK�Z�������}����O�r����v��
7�t�����H�	�&�������_+AEhhnόü��tZ��	�?/Y�fj�8Af1��%�g2�`dDQy�w�`g�ڦ1�+>�m̈́W[VȘT!9�p��pv��R�`�:(���%&�Y$ׁ�]xY�P��\������_��[��%K���#�ϙ��d��U*`ry�_�8#��%n�B��"~�Trb�[����cb�@1���ߪF/}�m�{!GRMg���搈��O���!q[p�˓�xh�0;c��t�x8��4q�]�5(����d�A�?_�gr��9H��Z��HVk:#S�n��i�	y��H9���Uy�Ji�Y�IP�\9B�:���>�~�����UcAԝ�$Su��>��zA�#
��S�kI*v8��E]pEٝI�%օL�$�Rjd��
�ґ�{��J����Zo��ֹ]����j�T$�\֔�N71��{�I�6�t$��zZH�M �(����vF(v5nܚD���b���Dҟ���0���S�-��O��|�M�Z(װـ[3$�ҽ�~����ʱ�טÜ\Ҕ����nac�ӓr{�A��vk���%3)�@�~$�X���k��n7�E�Ů���kp����ھ?�J�"��W���	.}�M)(�J�=��ͷ`�y_�<1ǠUw��Z8#M:��:�;fG#�d�b��g���xb��Lv�V@ƣ�5a�}�^��2y}���M�B�m;��F)����8#h4w�E*"�y����Tf4ԡR�ܤhI�20ܣ(��Շs���W��՚u�8���o .�C&�+g�����d��L.�'�NT�~��)r�SIX[L�dG!S�>@�����~4��
	ry�x�6�AYɗ�3�ˏ�k���k|w�@2�]�٨wЉ���s�} �����OYkY�d<��P����U���V7S��.!��N�����I�0��G�o%E���tU���R7�_���wچD*����-ܬ��T4Χ�!۠���ܗ��U�Jy���sHʷm�N�¨��p�5}��`�k<>k����*3��<e�����:��p\���:����̇х�"2�o~x���գsb��eR���3^�w�B�o�g�];J���s7՜Y����<�b/&�5G�V��휄#1�Yƅ����}���b� ��b��Ot��QyX�֤X�X����ϱ��uZ�t�]v_�P�����Y%Yq"�#�>���}�]���t�����#�a[�K��<����v?�"����4vſک�R�ۋb��]���3iČfE�'����1a���L�׋pX�/X��bn��ж�@�身n) "�ߴ�E����b-X��Ke0>}hR��1i�9�sz������	ѕ��޺=�����b��ԥ���§�=��J�}��#�>�BB?����lW��j����'�����d�M�+�K�Γ'�\d��<"}ɪp,zua�իy�:��9��V�l�`8A���Z]�I�tD��� ����W�#��,��� Cb*=�'i���:R3P��#HBMߩ��� Ĉ�_4
��)Ѿ-V�����BP=��ʌ� �,�����E6R��Y���P�u�Pp,�Ç�|.��a����64���5��-Ek�󴿌c�P ��ﶎe��s��à��*\�`�+�-�N�>H���i}qM�g�>�u�8��QF��)nL�O`�-	̈́%�'�f���4��ϻeJ�v�k�HX��Bc��cs�g�q�Ҹb�.L�S�a�6��,� ��KȽ+}���nb��ya4��QԻM����譤�e^�ͽy�~�s��^q�zB��#M&���tG��S>�y`(ˇ�(�B����<��_y��ns�V|n� ��Y���8�RJ~��Vb9�4�[�		�5pZya�S��g�#;w����d[����`=�{y�Qd�7�ދ�E��
�<�6=-�z<M/���+$C�=7�n�/�ct6c��W�	"����S���~�W���Y���YXz(o��BT+��q�Em��0p��ÌB�xY���^]��1OQ+�'��4�Jg���R�$o��xSK�p �7s'�,r�����ֹ�x���,��Ig"�v5W�b蝿_9H��}����^W�;�Ӿ�5�Y��1Nٝ��֦<ݡ]�zK�萃�zC�1�L򬥽D���8�״���E�쓜�~� 
�͝�6
oղ�.�#�@����T=��ִ��'��f�L�� ���oY1��Ǘ�?6��b���;Rm�V*g��	��$�K�j7;T]c�HW\�NЌծedm�ҀJ��6Ɗ�Ml���u��Jޫ��z�S��bǷ�m��|Ml��ɾs��{㙭/w����&(1ɐe��cq8�0-:�P�����ъ��4��,2Z��5��{Tr�~V8��vm�a�
�؜璚e� �mۙ���@*f�`�OK�%��'{��>Ent�5u2�0��ԡ�I�2�B�m��J�9ҭ�������Ì�5��u�WxPq�H)��)1���g�O'�,������!�%�ol���4�X��U�fgUr6����/���	m�pA��<���$����Iy�d�w�W��#}�4����:NW @�m�й�#�F�{���10��
s	Ű~����6є�)�i���x���P�����6�������E�|��ɚ�hWv;o�@CG!��]�k�[c�8?�L`�G1a��H�����F�C]I�m�x�h@��&���ş@X��;�C�7Cm[K�z��\oT����#6����/�Vx_�F��r�� a3wo3�v�!0���S��+�.���e�|DbG�5]؋�o��F�eٲH\{�!T)�%tr�Zѥ� �"�K�ey�	�5_��#���ep��0����/..��o���kٰF6O���7Op��B����>�.R����l ��y�v~��ڭ�wU�˟+�Ï(�0�����}��4˴�M��<��qt�+L���U&��@�[#&�jF��r�g���g|t䡖��6��Ɵ�ߊ3)A�������=�5�!Q�?O*��-��c>֚c�*G���k�Lq�z�;�M%=�g��a���y܍�����0/.^3�i�I>&J�}T�|c}vP@�e�Q�G5{�,K�0���F���y�Ǣ��b��k`�����p����Yu��:%��I�'��p�E�w��kV{�J�9�x�jhAY1�lb9���������>���J��nz+��$ ����siv�9��K��Q�
3iI��>���i��6�^Œo���uu�\W&{��r LA��g�����n|���t��ps�a{�QO�Eȡ��4�=��<ER�0/`44i��e�֘�թ��7����v�d���ٴ���z��s�2x��̒N��8KIo#;�pJD����wC�$I�zqa]��^��%"�}1M&�!r�Ya�gK����N(�U{���Z�MPe=h���3�QZ!J��syا�7�ct����gкm��ax�GX�����z/.�)�ahCG�^�祗`�SE���~P��KF>O��+�</u˯N2��3Z�̴�+�դ;\��L����Il%�w�����{���oC3��/"§���S=�}�AQ�����n=���c�ҏr���Z�A<˳І�M*[E�gH��փ��Q�H��(���|�RaH���]eR���Ԃ^��Ήg��Ny�8�6R$�D�3*%N��F.��57�JQ>r�0i�M7	���@��2ox�<[&A�Jϛ�a3�7���	��Ҧ%�}�!��$�"{���������dN�/��`:����P�����hDW�?�{��
L�	mK�.�~�"~c/�&A�f?p������b#��3g��DSk�M<_w0��ߙ��Q�'K�C�rzmE���P�HQ��9������K\�Yr(�~���O����6$�#nԺ���)��B��;J��uc@�q6Sn$c1�>���?V����e1�)��>8��d����J�� �
n}��kcb�ܛ�*/[). �+�R_���~�I0L�3?�)�3��s������J��+���]ܴ�+`�nt����@u�&5�QD�58	!�x޴\�c�))g�#1V����RڗAM�V?�R�^���6�=�����i��)���n�j�P�o���[���1<3�"�L�"�>J��ë���ޚ��0��}ܖN9�8q�`>j?9.�Z�[*%�����?�T����+T�1�7��\31�r�̔h^�� h��$�">�A�X��(�K�6�2+����� g���,Ep$���uh*W{��H�~���d$r�<RˤJ�%��z���d�;
t�黃�0�v��akh���s��w���*1��xB�r83�x�S�;#̏�7:��&�l�6d�O�ǿ��}��L��C�b�V2�Ni
���-�˘�Hն��3:n;8�$�/	wHCur���O A�e�5X/%�8,B���o�����oTK��H���
#%����WcL���bz�Nb¥,���Z@�"���>�Op�璙e����ת^��D�U���e�����������|�,{�(��m�	AY=��P޲n�}��nG�SD����t��%5m:���>��m��,6�~H�={�~)J%~�撖�KP���5�v|��e�x����|*�D�:)T n��[e> ����.X�G˅��k������״U-�L,m6�%MU*Л�A6
>f�'�Ԫ/Pv`확a�ҋ�VRC�P�ߛ��GxdE���/8^A��ўu�I��h.Tu�f�R$xt���u��h�ʮx��'��I�`�.*<f������m��Nj�3g"��e�+`�Ư���Q����a��@Ù�����c�Ѵ�}{Ӄ�M�|��A�<:�4\�0�RR��<~L����I|����}��h?y��p��i��f����v���0���|�ׄ�zȧ�x�6�k�y'�'n�������k����;��xw�@]��2��9��gJN�cOhۀd���[x����"i�����r�6���4�~ԴŮ�U�Y�+~}�{��o����s��6�$����Z�Ѩ�*��w�Q�ĥ俵��#��0�}�֠bt��@/�&b�|d�ܸ�.��e��t���A@
"�a:*��ΐ@w���g�4PY��eJ�PoųTtU�J������@&����	j���.�٥��?�������F�"&�XOS:��������;a�ёsF���f�=`�`�p1�P�)�ib�9 ��F������c�'*{l!KEK7�m
o[<�&S�n�^��y+YĠ�h�ͩ,
�v�����g4I��W�����n��w��}�v�.-A���-<l~wQbW�`Xgԁ3W��t��� ��Űk[fFje~���䅍�lRpP�'��_CM�=�Dp���u����r��y�������C�:("����͘���g��=��)��S���Z����.���a%�@�s%_�~5UW�ӜЛ0�H��N(e�:�j8sLb����g�Ըn!��k�?�?��Xo�=nvAb�<����x�=���L��V-�� ^zd�9u�}��B��at$ϐ������1_���#�ei�H5qA�%�����o��wD��8����jݘ��Fw���N�P�G
�٠��1%�{�c�c@X'����w?O6ڭ�\@�N������p7K��Jp �J�,�k<��������� �XHom��[$��9�D��6�c+V}������ښ�F�%������˿(pe�m�*����)���OI͸���)l�r�&�NKbs�d�"T�eP�E#�eph��'��)Ø�^ XT���\��B^��VZt)<mW���N{:��}���nU�!�7�D`��)�CZ�,n����!����qڒ:����)�ԏ�����nJ��TT��)4�B�\���0$�U�p�=��c�vP��_ ی���nX�pL<��joڽ2�������'h9g��2NV����?�i׫>�$U��v��3/�}�Z�0��-�#
��Dwz�o 
���廜�M2x���2������㮍�%��8���^�)>B�%�T�����RU&�J�IYb8>�����Վ���<��];��E$����g⣺J]M�� �M��&�T�F�wZO�������6�W����4��k��p�ˉ�x�i�>Љ�K�I���<͘h���*Ml�Ph�h���0��|0~�7�E|����(�ܓ:^υ�	}W-�f����z�5��iKf���k���Öo����-����mh� ����&6J��БJG��X��r�^v��
BI*�SV��j��5E���L�[�o�Y�������X@��̸��;�"�N���أY.�io�o���=?�^����5�OH�}U�_F�(�ms��
�1��ey��8;�2�)P�\p�x,|�������P��I�˄k��:dtXn%�,�$y.�0]o7r�4WO`�Rq����£��m9UT��Ŏ�w[TZU,���E�zN%ku���+��l<d��c_���V}UX�(�O�URl���~�G����xs�`5s�S�����s�_f��R�\eH�m��	m�/ٛ�ϝ��z��r�w��)���k�8���?�'�:��DM|"W �TȚ�cZ;���w�\B�{�[���䷃�K��ڐ]���q`bW����Z���Ġ�֮�.�)����#�����^��V��s��Z���f���$�9��V�i���YW�3��hɚ�	���Ck�M��T�����O�^R8|̍eI s'���Iɟ�\��ЛJ�����Y�(GO���	y���9s�ɬ���p=�b�Z�� 5zy��է��	��癟�VJ8d��(�&/�aUmE�)�c�����EZ�ܾd�V�T�iM���g�c�CE�Kp��'=C ��x�c��*�Vm\ۙ�)��R�t�� �2С1�K��6��p(Lv�o>�s4��[&��p״N�K��M�bn���'P\ͼ���K��͈��� /�z�o�$FNe�����j31/`P�E���:�FWc/#"���E���n����u��JE>&#iK�-6�LJ�T�ҋB�
t]x���$��4$q�xb���M�G��ӱ����?�Ƴ�fa�;u���w�����`�X�uZ��'��N�φ٤�Փ���16��D1���Q����gG��N/g��ܨ����n�F���+�UL�1����10�Y#n����f�@�`2�a4C�x���j��G���D���Fc�s� ��ln�Lb,keW�]`�	(P+����@���H:�>_QWc�?D�T`�H�%aGU��ю-ڂ��mK�lS�/�غ5�2��D��&T.\}j�F�y=g�A��8[QG�F�ʓc�������	 �<�n/H�Y��DO�L�z;�ݞ[�$0���߁���W:��0?��>Sb�t�v�Qr��%a3!������`�������x��6���!��c`�<=�}��ib\n�͂i�ۢ���~���i5�!^�q��c�8�	�=b�w�h��ɛ�=FPQ?V޻��+�Z�����`t �,i�	���{s��h�b#zK~�m�t|�!ƅ(����61�h����t~/n�&HV�;;U!H��>A��_��~|�/���h���q?�	
)?��GA��� P�;��;`�4���eFY���g�Q_İVZ��b5�2BMٶy PV:�+�BŹ{��2r�<'�$����	T�'�L�ٓ�5=��?��0������Gg�L�Doz*cqa2p9p&4]�z@�B��� `�ڰ� �,mMv��߬���	���k˴">��(��Rfß�ѹ�B��ݒ��E�Ң�CO��f�u(�ީX�)k��$����4%Q��Ý00�����*������X�%�pq�-
?��K����]��Dv�Q���TM�!�W� @\D$,����֖�ϳF�m+��T�p^���5�G�Ԟ�o{�k����>� 3N�y��E8CXu���lwU�oN	����z���)j�!�rZT<-.�����I�m�:ۚ��T�%r.��>�mu1�V���{x����n�a� W< ��_��*c}C#��F���7����G���L
�.x/c�5'����BOˇ�ei���3�yu��~���v����<�MX��&��n��ګ.np���[�
�N�[�T�Sxc�����3��8jvom�{_�m��Mbo��D �#�q�F.3�I]��4̯D'��xR)��ԋ@��`�C"��X:��ݪ���ʮZK��kj�|*SEC��7�����i��U�`}��z�D&�O�C���t��e��XA�`��(�+�H�ٳ�0�`j�ۜ�r0l��6rW|�dC,Omt��E0��X��7��x�E��/��H7��!"�j�I���E�w�u�E�"�I`'�*!]�OW�#������З�>�_̫�S@Lv#a{��kCj_�8g?ں�N��b���tmB�Yŏ��H���&�@IռX��E.i����!��pI���i�#� Qƨ$!���H<��K�ʪ��������v�]��Y����qo-C���(�Hp{���ψFO� �o�)ɾ42s��v��̟W�����i�DjJj]1�?�p�����3�pgɌ,\��b��Գ�qϔ�����y .�|FY�� ��Us?S���5,��V�f*�Yx>W��d�e��$�G,h�8h�U�	_!�`[��H��;�������1�<���|L�����>�iyV������5�1�PTmTF�^�n,�,�A��V_4����e�]�gk2%۠����=�3�*��ѷ��[��Y�&����(-[�!����b+��'���� L�;v1���yY["iK�&˼�Hfn9��ݽX�m<W7g��a���ΐFV�����2�H���hg �khe=��M*K�S��l�\eM=8�3����(�kDJ�jK$���pSRw7D����፪���I�e�Z�P�o��k��9�I�����V��Ŀ"ݴU}d�0	�uq��^�C&t8���ѯ�sةn`����
�n.M�ĘQQ�	q��Ǽ�쾱D��{1B��NK���,�E��Hx���Wa�d6/~?QX���c8��AT�6"ж��K�=�T�p�L@�;r���ӳ���͸�M���R�e�<�R}S��6ˣױm�71Z5$����[��/�V-��O�~,�Ђ����7��NB��� ��4�}eVc��G��]�
�8�6��x��s���P�/ѩ�bW:�,qqZ%�EG����� ��r�mk�H��٫&� ʕAsy$��?bܘ����vkFs3��X��K[��*N����O��Tc����S^�'�1l0:/�?�Pީ��7N+�Œhu6������@QQLݘ�2���{E��2n��[6��S����c�2����Y��%+6�[�g!�-GU%�E�4�A�z������y�p*��aS@��q�&Is}(��e�"���T���Jmz�Y��l�oƲ�Ҝ*� OL��
(/6�Rt�e�(4F�����~��ǝ���t}h��t�B��a�.�)/�W��"L�ޞBFը�������`�hx�Six�n����v%А�[D���VB��pd�s���ĂW��:"���o�cz7u�i8[3'<*JTό�m�i;��W����H��lU�E��J�)M�+�)W���m��pн/؋��&�r�F�z���@���Mi�ʗ,�ᦢ
U0bǇ�0�qtx[���E'۪R�EY���;��W�g(���67��H9-�D�_E�⋩3&���6Z̎ā��j��r�9� 7C����,�l%ծIٙ2|���H�Ru���)�)��nYw(A������S\�����h�|��#k驗�Xf|#E 4��1Q��[���P���C��ȁ���J4�kP9�z�����d��J)__
�q��<�Q�U6��뺒��Rȁ&�<�N�?
n�w^%RӤ�ln-U�I���<Ζ��pR�*��+�1�v�N7��5���n�^q4� �~Pg�%�>BKM}�qUպ��9١��i��e��&�J{��	��Įpt�D��eZdY�@�����sj��%5k�$U�\rnj\Es��`��Q�a�(��PT��ٗs�읞1XĈx��W�p�Tfߵ��zH�)h{�n���̻E�MoF����3�3g`bHxk{��m�D������Wg�!V�Y�|�`/p���ѷ����ŗ�$��`��K?�ni��+�*u����_� d�����@�J2$E_~��H�i����H����@��Ϟi����~��|���(xMP���k�ũ���4M����t���N�3"��yf��sĞ"�,�,�pcc��˝|}��<������s�<�s�VT�����g����۝�E#DQ ��hL�#L�f�s
�Q���)H(&�_E�-�����My�YU[y���Ғ�����.�?,��O����=�"�،��[3����������[��"(�[�����I:ԇ�v�B=QC�
^�Ԟ�u�A۴bX��R[N?Gv{� ��D�M"i;z��r���Wi:L�L�	*�GVgE]�2����R�^�H�H��@��H0�}	�Eh�wf�%�X�NuHyE�z�d���}Jn���V�q��x���{�_h�q��3����[rj��F�mH���� ���SCi��̨;F
���`�(�9��]�%Q�	�t�98�����������c���+Yq���tdVa$�����.קE�,-��S�y��&n�g���f����D�X�BU�_�ȯ?&���z���_���DFN �8
4ճ�����j�h���u��L6�*���X�C�S�|E���뼒@`g����F���WX��g����G�|QL�j��'뗖��,�(^{�b	M�]`(qG(����&V�L]1Fp]�+���>KUaxx����^��{,�3��Þ@t����9�^n ^t�a����+�Xɷ5A����	�S����p�n���'�g��@���t8�E���x�WC\��V�� �`xL@J��[�p���g��QW�?�/U$��w?�c���4Vl��YV�rO��f�[�J�n�U���V��_���1�����O�����MC`��haJ�q�Mv@�F�ڨ�^Sp��Xaw�
xT�$lȓ{�L��ݗ�g�E&��������C�70<��
�e��4j�7���8Ec/<��>��ܤ��C�Wl�;,��v|V2 4:���8ο��ތ�l��r��\갊�=�uU_�̉�J�L�9���4��~�)ty�Bu5F�%�:�}�;|��b�uėF^&��w��5�]%~���9��un����#@���x���N6|�I߹�7�]e����e�C}�ĸv4�|
z�ٌF� ���
��O��+���,��coZ���l�Ǟx2�>82%��;.G?Z�#f���p	1��F��X��D���ą�@�a�4۽ךV�7�԰iGz�� ��_��{K�~�Rd=�Q�]�>�9��,$���-�#�]�,��B��Q���gn��bE��ޘ>���q��dJ*f�l�v��5��$�' -�ֈ�u��7puTm՚&/��a��p��ϡ�����y��ˊ1e�����o��$r(:'����!A,�ke|����uK������Իi-���B�f�w@T|����iZ�W|0I ��$ِ�/�Yo8�ŀ�F<zl?h-�%/���L���a��$茎��^��ׅ�����o"�AX�,��Ӽ�I�kZ���mͶ����^��z����� 	k쪭���rc-@%g�u!�;t:��/(���Uq �,8Z��P�6A��'3�����_C�6X�<(�؏�����q?�MἝ��jE����WڑW���ZmXi���@ H��ڒ���9.k�4���y��kjd*KÛ����i�k��M�ja���_��{t�nǄh�8T�3�%r�LP�P����΅�����S��Z�hj^�*V<W0��lXF��ce����x�싑���(��a?sՃC��jF�� ��T�ӥ�l/��d!���*-���d0 I"U �����W�Fg�}E�Ƴ�:�W�w):���M��s�ś8���5Ey��w�t[|��YZ9+U�d�������8�^���qNfL�_WM�~��Dgޓ��le����3�Oy�d����^��ʉ3���k�D[L�]�Qd�[%s����	;��0�k� K\'��>󶌍n�S	�d��{O�<��d34E�g>����$�V���2�V�^��H�ǵ7�\RV�k�m&����w�k8�����`�/W3i+�,�!�f�iy��
�f��:���	]�Vd��R
�X;%�}�vh f����>���@|E���΀���e��B���}d<��d
H����H���+q��=�G���Io^�L�4���zUy�-\T�������tg�г==O�Ȩ+[��o�[�0;m�A�,���oI�H�F��F�o���?�M��2�G�)a�5�������������+�rt�L4�؉�G� LGM߰��]m�ȯ�Y"�|����6p�'�"m����e���-"C� F�w#�J��$�䵒�q>S������.I-J�QJ6��,���o���J��~�b���[�!�ӱ�t��Q#��p�X�د����.�xբ�!ע��-U0�j�m2{K���E��aL�<�}I;���<TY�c')�ht��z��|�%�a��3�0#�F�R3" �	,ȋ/٨>z�Jc��]�ճ�3���el�k�������Z&2�@P�➨���Ʀq�ι͘j���z�v]�E��`��i�J��ͧ����v�$T�p��{A����εϨ�ɨJ�7��J\� zB��(�Av��C�R��
&�_�AXR�⩍�P�V�%�x�k��i>���1�B�Z*o~�-jb)��S>	JH-��_C�k�%IǗ��+ƾ���<�ڊ��AК��X�s+]jjfʶWGy����5!+��꿛����c��̋�e#���V8h�ΕiQ2$LLFv��y����# �lSz�*�������sL:%�P���_���Ա__)V" ��I��kL~�+[�I���l�]
m�u��fR<��Q����q(mx Zb J�4�^Ri��Sho\�	�kt|�������?�b�2��P|���l�G5�GDF,�U�[��K�m̤(Q�8���=�R�@���ƈ8�sG�!]ů�}�񉙌V�3�g(��9{O�_�����rj�*�@���q��5�=J���zA�j������]��K,�t����V���,���Ӓ⌻�}��O���?�JFn*U-�2u�
�b��l���!E�Vj��b��*v}�[=����:|��W��4��3��4�S�	�jG�q�r"3�����Q"�]��\(v�U���c�;� `��y2��[+����g�S�hKmѨ�#v$px�h�p�W`y����f�A��4�� au����%sE���x����q�=.+��O���%�Xё��M�;ך��
��Ը���	PB)��a[�о����A;�j�[(u]�r{�#�^�7�A��DE|+#��V���)���o�'�� G����t�aÜ��L���<�h�3��;T���5CԚ��F!�+-	�$azT�������N�$�����x��F��0˱�3A�����ɯp���!ݶuL��a��;�=�,#���$@L��3���#�y��<�1)�%��,���L���nEaE"�,�Վ����@Ȳ��"���l�����w4ݪ����r����\b��ƛ�c��
�dk]��}��_�CY|��;��s�-
"���֦��9b��N��	�I�.f/ �����M�d�^�9^��o��]��V�A�%(�~X��WSq�n��l����Pm;Zt��p�q?Ÿq�\�\w6��Sm�y�]��Xc ��{�v!�u�X7���` `��L����S��',(���i�~tW%"�٢,Yq/g�X���"%����:<|�5�HCK�����k]E|c)B�5��!���K�>�*��Ba\�g�^A���C�t�>[S��ʵpZHI���ќ���̟�/T�$U&]pT.�c�s��5ˬ���X�N�|��Ö`3osb�1.�1V���D7�(�H+��催'x�*5�vh�O�V�f�t͔��ٟV�� �3`ï[=9�K��3H��!�"���F����o�{֏����.�y�U�!T�M��pF����C)xmT��r��-�>��5��}�.���s;A�!�1�_�l�h�ybe[�Ge�'R��By� DCt��\fvJ�~�����5���d?r�=���!������@W?d�K}
�1���#���4�	Ṿ�y��*О��T�FLV��
Uϩ�x�
mW>_sy&��!����rV%�"��������N�rN3�t
���3&��4S>��ȉ��{�k��fǂ���8���lRՔ�	ﲾ���.��lۜ� BZ����-�(�T����c�(�2��cVot�t�^����%�;����M��ݓ�8�i��N 9d�l��2� `��ZA����TB�&FDdE@�{��p���Qy�.i��0!'�5�LgQ�OX֎8t����tC�XcmW�U�����.E0 ;�7:�
�+t����'��H�s�Z��N_����=S�l�G��\���8��#a�7ٝ[ &~��$_t�­g�1�@D#���Y�q	��F�+�0�L =�}��\�hB�ﰝSq�&�2c!6�	����9����I��(sV���vªib���4��䲦��h,W�Y�x������r6��7���] �j�B��8Ŧ{�[����m�������`�Ηx��)Iyw35�S��+����3iy^�B�Xj��]GfG�K<a�xc�3`+C��<�S��������(��q��$�߉mF��N�j����$�* iƕ��2m���@,�[�񌫝J���.|�,��CK�� ��������j3��>�Pf�ۉ|a<J=1���`� ]W>b��^��MŴ�ڪ٨����;��.aD�#�g҃��7�i�����2�^#%s�V-�81z��5l1���uQx5�H���mu{���J�<}�= ����A�����D�)A(7�p��pE���7>��
_�0�b蒮"V.���5.�o��J>I5DB&{�Ģ�i�n���Nn�w<׽ב9�H�"�� &>�RK3��X9	��_H�K>�W�.�i�Z�QP~2}7Ĵ���w�ԇ%��z@��(��8&��r+����:��y�v3'�-F��0�ʆ�Us�v0�iF�}:�V~Yd>�Y<� ��[��зY?�U�󄝲��h�W��u�X���|֤�b�I��9,Ỷ��ǆ4�W����� F���#��95��>������mb���U[Yc�`�����T2w��4�=.������F�ZR߻ZUx�zX�$�����x5�"��=�,�p.���C{"�����T`#8z˱�#�t'�����U�\�φ�-�ς|�GfWA�	�c_k	1����J��UE*}U�Iqa�	1�i����a��T���"�$���t����l�h���n�D�i�Dr�(���ڠmx=���H������o�C��B6`�x��hǜ�>�!�3n�@�q���@'W)�-�ð�"K�y;�%\ø�t�r��߷�}~���D8Fw�=�v��l�Āc�g�u]� �$�������[��JA!���9+U(�3��m|]�`_�$��f/� ��!��` k����qԾ|����~�(���j�����ՐQߔ�2C?�����j�Ą�F9���٥1�0
_��FXK1���7VH���ݯ}�nsbؿ픜-ݘ���|��>ƟH���\ۭ�K!�c���2j]?���8�ԝf��rɠl61�&�^<�v�����@!��7�G�!�}P@�2iv ��(�~=��p�3���
���\~�v LRf�<D>۔Z�<��i�nw�8t7|j,3�p�
�|����"����6�����s(����!"��;�$	�O���#j�XR�6��\��]�ÛR�X\�6�Γ�TF������$>c��e�P,�ʎp�wP�u��;G��}qd,nX���"���8ʹ���¾Ӏ\1��1��WR�n�b�~:�rL�F����R�@�7p�����������ŉ�~b�E7��D�Z,�L�vt(j3�T-��	�ʽG�#��re�}��:���F)H
�����?IusC���I-{��DA�jx�1�<Uu}�-V�i�\hW.R�Z�&��)��D��p���8�ӛ�6����-ݟ[1�RA�o��a����$W1d���L"��1YԁL&(?I�,]Xw�m�o.�<C��rG�g�F�d�H:�uA|K���&�R�;�3�*E{9h��}w�М�o���N��һ�H�0q�L�'�SP�������g���X�|�h	�l2/ULz0�� ���4��oc��$�@cT��Oh'y���:�`i��j�Q}T'�h�!���r���dv)-�� 3G��	�0��s�ˏL��sHѩE!��6L(��n��>(T�߉�������6e���;cDkI[���㺮Lw��C�#ɢp�%'��7���Cu��Z?��ބƷA��!l���}v���TW7k=���~Z�D��.@"�r=���9�I�vT ���e���藘�b�@�**��p]������.�<�L����p �6�%�/���g��D����[AE#��l���eg,�\(V��n��K�<8D��q�P�x�ʟI��֩��J�뻰�d�yƨB�L��շ�� Q�O˺�I�h�,#_r�p��}:���1rJ!X�$h�ƃ�!_�v�wҙ!�F%:Y�}o[��(mF��M�ځz���m���62�i�x	�74hП�����K?�>���嗢�?L�ϕP`�߽�p��Pv�`x�ܭd.e(
��A�sQ?���i�/}[�XN`�;/�M$3��'�<E	�� ��ۼ�����L$��?�p�����=k-%@��r㲍Uο'O�'������+r�"b��[�x��`�b<�H�����u/+S�'�ޢ�e��`M���8�IKR�� ��߿�`��{��ġ�6�uؠwQ������F1A8��AJ�c=?��O{Nwhվ/��u7ӿ��%	q\��n�=�#�K��-��{/ �db�g���U`�H��!"A��d��Z㷗�q��{��@���R����ƭ��j�)��,�6m�Ʊm��+K݀Nw�A��0���r�T���7�w+�]��0*"[�7*�pBM��0�*Q��Q����и뷰�� i �Z��,+*e�g�9�� D�a9.�_3��j�M�,y�J��06d:̭���*�^�(.?�*�֦�x88��3:Lp�#��%َ��
��zK$C2z���Nao�mLG�]�-Ruj��I���l?eE1�O��TZl�ֹ��ٺ&<U��������z�K���/��0+�3�'��H��>L�.������w2s�qbG�֮i�@�S�:&�����7�o}�˹8X�P��2�j��aQw�#;� 
+dQ�]��J_E��6R�b�:�����WjS�=�$I0}uk�#���>4͞���F�ek����}�o�M?�d��+Ȇd}��	@�W΍���A���3�M�ì�{5Aq���hm�7� �r�"O��gܬp0$ڗ>��YH�s�O?P�T!MB3��.W���އ2��T�­_	��tr�����eU|oNN\��hu�0u�\�s��kJ_ԏ\Y�{��)�.�:$�ў���X�lZD���cי2\���i�zˁ�����e�������yYH�7��xE���Xv%
q��-��ة���[O�G��!&�	uH҄- ��b2�!�hC����7�������CJj�������U^χ��v����U�'LK�C�Xc-5��c��2��q�>�)-�`4�=�dX�dG��#�R��
L�xX�/��"�c��hG���\�ص���&VF=ГTa�����U.�M�RG��R��Z�UlE�W��h|y�v�i	�y���A���p;����`�d�|�{��]��£]\��y_f/��k:��}�ץ��駪��	��Ef�L��-�.6w�Y#�!e���[�8_��-�d�l�����ŭH���`�g���~�<��󬢝r�1�!ǟ*�͆8 �aټ�x��C���VԽ�9�zk��\��m��6[Rk����X?B���g��i{Vζ=��h٫8s��r�J�\so�F0��V�a�P3aVW?�R����R�T.��(VM�W���R�����R�ǲw3����Fv���Dgpߊ�;���0����\^M?��F�G�Zt$�<�,��t�����b�^�՝;�������l�J�������Z�5�O��7�ҹ�V~��8�MF�Y���9+mL��&XmI�j����Nj�B���u���k�R��h:��D�9�<E?�5����@"�]B���d��<҈ ������+�Y���.�5pO�|�08ynS)�lR��@���[x�<+��Km�-]��w������狕���#" 4'Ҟ�q!��,�s�A�^��gˤu~�V�^�������.P�F�F�C���q����%�^q!�;XY]��E�n�I�$�׹Km��'��������*c�d����Iռ#�р�w���.7~�&P}�$b�yx��x�%�6�%��]<�H���D"��_*�jb<
j�#ٵ�D���C��Q�$�ʤ���KV|?�%cH�|��DO��/���dLwhظN3	�����YM�Dk�tK�f{���gSJ��f�{��}�gu��:��6�3�+,'��(�&c��Uu\g=޹����?`rh��'��W�_�O٩sMoO�@�&����[S���a���)8)	��Gh�2au��,�"ϻ�������7��)��a#X&�̛U�ꒉǦ�1���j�O���;�|�5�)��(�� ��z�.��+���<�>�� ���ת�	!W���6��1�!�~�G��T��� �C�L���6��Dk[���~�%*����S4Y�k�6`�'�[2�w�)ѹB�_�zd�qwX�Wt�$�8�ʫ��ȑ���SJ|8����ʫ �"ih��r��(񒀂	LB�qo����D��<r�A�����]���	�<���kߖ�cH��KuYG�a��Z @����]読Zߓ���;�[_��>a�g;5Yvw�1��6��rX2	��Rݦ+�xOZ�j�%��aՍ�mgj:����̝�s�N w
U�o0x�����{mE���؟ �TO��?2�#��zkqm���%�%���Hڪ�yDxi[ ���Rb�g�K��L�j�o�'���F��W�{�e��X�9�3��+��gv��r�$ };�c�Y�^%Q'�M�k��Ń������i�G�O�O�yP2���𮨀MZ�7�*;7���c)Հ)2Ba��� ��x�	x�V��zP<K`��5͚/�UȾ9�)��J�%��7>�����]�nl�p�һW�� �������i�<��Fx=�?��=`�g�b����sh��)�0���H��(���������ϙ�I�S"0^O�9]75�8���R�wh�-���J��CHx��t��k
�^ j���^�Pl�w�ѣ#O/h��w��/��[3&�L�y�
�屨i%O�(x���$�t}�h{��Z�'�᧴h4�o\/0=Pn��0�M<8�4}V�A�Zuh���l�wի�O!vp�?��0i��qXK���|�8���Έ5�W�wWwdn>�P@�P|o��R�5g���`��L��b8V|��G��������N��!HÙħ�N�71'hZ$Qt"�OI����� O��x��S���»�,�e+Y����-{�c���uw ����@^����h��-���,
cإ�S�j�?���Y�"*Ց�XL4�/�#�����z��*�kE���>}J�ҹ�����	2�op�A�/�_}.�я:j���=}9�-x�дQ�®k���m��Ոӎz]�9���o��+��"���A+8��#U]"UJ�z����&�8-T7��q�Z�	
F��e����O�LLXY���|o���m��a��N�[I��X�C͡����S8�Hxa��z�̄
�Ug��C��O�����
pc�N��܏���y��+ec��zZ�~�-P�Y���+���ëX-h�&��B���ROq�0g��4�P	�7��Q���j~�#�؎QG,��.\�ɚ�ҵ
:�A����&�x��^;����7�g+p����3�F���u��O�0��	V�A�_��^geV�K��m��<��!�8B�M�x�L�I9��R7���Y|pEZ��$��@���g}�J��$�8w#�}�ld}�'�����fH�t
��~�R�^0����A�.f���^g��p�A~5�^	&}^���#=Ȣ3��D��΄��)�R�X�fĺ�?)x5��e�bZ^e^���{MJ���-�m��d�$j�f�T��^�i�!E�[C����5�/�`�:��_����Kf1k^�m ��
	�E<�ԁ��%q�HEY�X�����SX9�d�f{�����3(C� ���1��unI 0}����/�D�x�������ӈ1֎���
t#��/?Q�1���༐ �}��-*;o�}��Qz�xn�mނ>���ye��&T�g�-ʩ���[�H%2��^rR�q��ҜD�Zas ��[Χ�����KF������@ɹ������������Pu�_�?�P����+h��9�	6A2����o���*m.WUN!y����R�?9�����d�X����������Sf�v�h��Q�Z��ːaRv^#�0�齦 )�N�{@�_b���9�J�ǋl1�pɨb?Q���a����َ��c������"�0���!��`�vX���r	1����}�j����vx[�8�и��#���>d��\��j��E��ؼ��[nV$Y\b��<B�*�㉗JNY�5��f�����9��<�)��L��z�ԇ�K�G�Rۑ�	���������hK��g�Wj1���^���h��F%�nQ�w'�,�<�c��3<�}���F!�كG���?�����ݷ3�;���껈5f����_�12�_���Сh�zu0�-'�����p����uc�q����c.����P�k<XR��K�"WK�wZtF��<%�H����*U �k�5U�����Z�٘��	9c��@x�k�q@HmN���l��\�ǳ�X�+o�d���ET��������t��O���#H�Fn�����#�_��+�G��_�6H�Y$\@^`�ztC��.���eK켢�\RX���')�,Sr���ʋ�n��R�$���9�z��0� q���	�(���78�@�4�g�)"��S��"���l����5~��RY�9٩ބ��(�C^l�`����.�ӑ	�����^=[��ZsbVd��Ѣ=�������B]���6D8M��#�r\)�*�%#�Y���0��쓎\���%��J��ZJ�g���Ğ���I6��N�����{��#�
΅�J��A����p�a=�w�t��5E��mB���jD"$ɃF�	僼�#���:�د���n���ˍ����D�[Zuɪ��Ԡ8�-�zI��:-]�&��y�X)����n ��F�	W��I��,�('�Wv$z��8_MPA�<��뿻}���H�EjeU�3�g�$�Π���<'�$ǹ��[��W��_�h^*~��3۽��9T��9~���A��5J�Du�0T��H�T��"3J�=��8%R�~�b�ĥ�h�8�<1�Jfn*�z�Fq�ڸՁ"RX��N�w�6L
#L*�D�XtO��4��,sbV��}�>2;֒�*��$L�E�*�0��ob<�\��5���Q��52x�E�V޳&B�Qg��	���G���P)@���9igݛ����$���������8�`j�e�ܘ�CjYƴ�k���ܙ�0�^!f�)�DG�<>����Bmz��� ��L�m��.O(�G�[����F�ϸ�TF��y|��7Е
�0\�؛ L�0�� %S�������ULw��˧+[���� D��0{�gU��/?�̍�-gA��/���u�/�-e5�M6�IA�����ס�dH��Q��h��үG{��T�"�H&��mum�?BZS"�6�FE����h%�(�wh+��kN��}��h��nN����$����z,=�M����i��Lz?��PL�Q��1ȿNtY�Yy�����p����4qGIߜMN�ϖ�;V|�ky����������׍'�u����}���-���jf73�����(ka?�TY(�ϵ��{D��eB��K�<]yz����0���VKI�.X]��ML;¦ �Y��!W� ��L������#d�T�V���i̧D��q0s�H�A# ;PR�w"Kq���b�z�7Y������~F�D*P+�L\�MS��7�����`XS��"�Bz@����m�����2�,��H^��9F�/fbn3���u���b��"p���$�/��G�n+�
ٌlE΅���]�M�<e�X�{�T�J�(���b9��c77PR�>�XF��/3��V�X� �1W���V��f��t�����t�:�)�9�B����s��7�q���dB³E@�S�1!`?��co��
K:���F��j$��+�
����Jݤpu$������3L1��蟺����2�9�Z0�_�@Lٔ��	ޤ��k�7�<b�bnDS3B�ԢR͹��0E��,/>N�ܴ��wp��s9��?@���B��;չ�*�Ƥ�����-�^r��q��V�2�׹���5��#������=�}�)������?m�HSI�{��S�}��?��N��������g�b�;�$h��|}��Pl�	�Yr�D���w>L_��N6yH�֊+b����I�q��$����1Y'\�G#;[(Zn��k�{iv���^e� �託8i�̋����< ,8I��6>��ҴXo�,])-�fU���?x��  ��Z"�O��}`�˿¿�R�h3p"��9Kޓ�i�	�ܝBMDy�s����i��2�40�m(�J��B����PeYeҼ�,�a)_ѹ��:<s+ma$j|ؗD��h����	����4�u��IC&�5��-�Fy��s�~�+� "����~*�T^�� �hz�Smv	�X�*%I��e�f҄������ҁ4��U5\��m��-�fq�^[���ǀd��\:Q���ke����;�@b���6�f�w=��fF�NW$��w��� �䴟�	'A�U2H�W�#�e�Dq���(|�[v/V�9�aB�H�6w��a���	� �ҭ��.m9�p����x.H����U�y�)mcf/.H�+�p�nN�J�Wߴ�v����DE1f�7u|Pє�+�� %Շ��]���ldUl{
G����$26�WJ��m��&t\Z��pohkf�������p�3� o���
���l���㙢��@r��R�pa6t���G@�p�z� �$�I���6�@�Gh�-�������)���L'��ؓ��B�@E�ع;i�;F��4-l�>LFղ�HR��T_r�� �1u��׼�Ȓ|	����� o��_0��}}�/]"�v����_�nt�1�8���49����pI
a�H�Z���#�/vj\�r'>�_7�iP������24��m�|O�7`$�y�=�l�S�T©��yr_A����(�J�z���>��A���@�M�u^g��\��j^�Ei���T+g��Qw�S!�L�U�����Em�ew'��JY����Ll��o�d������^�
Z��yܞEa�o�����!��B���=LL���P�Aw��Ӻ-)�QSw���wWP�c�/���1�{-R!ù@����.6v'AJ�=�sj�5�{WR���6��'��'[��|_�c��	��-\yC�"����q#�f
P�it�Q��T{�[�}N@W�b�{l�}��\�Wd�!8*bˮ�kg�PKp��`�������Y�v�N��_~��X�A)�*����I����k�Z��Ͼ���re4���Y�R��3��wя^6�c��� [m%@�(n;��	r�����ߘ��+�������\�����N��0G�ÒL��V�v��l�D����B#޾b!��ye[�*e���ӽ������DΡ�G�yp����@�T]���bݡߒ�[f�N���GJ��`��ӫ�j�[o��8�;x"��Y�Fh�WG��&��T>���8�=}�=k;	�u�	z���q�JЌRK�b�j�ȶ:������;����f��4��5�-�Y}"В�V�oq4��`7
0~�=8LI��b�H�w!��ge]?T�uqA���Ꙧr �������Ӿy8$ڦ�^�.�)�%��4^����	��@0b�~������'	,W�؟6g2G�M����cW��c�+�︹Z�`��L�&�lo��hֹZHu���0�B<�m�EjY`��i-���� ��,eV|k���'R�ɮ��+=���p��i�SfIq�u�.X�,vcy��4Xyn�5_޶Q�դ97>UݻXz��{ϣh$:����'�Ld�,n�w��LR�_��8?�4���#^:Gt���'B�E�u�V���,�8��0����l�\��\e�&k�I޳N	�T��,��(ް[R)w�����x��]Ka$�F���e����y�}&�@�)�����yM(2lu��p/�H�T�ͩFHC0�(y��T!�S^��A�ߘ4�H1�X�}�P��K�xb��3ә�?�w���A�:w��¾��-�]�KX}��ɓ���Tf�Y$&�6=䂾t ���"5Ð���QO�$� J�g���y6���pH-�C( ���J�nZ"`�|C���B2�KNy�<^����BQA�<zs��ĕ�{�Λ����y���k%�3������.�ɟ6�ȓ!!}��]6�s��p������	2h�����������Z~8���������ROO�0P3���yݪ>3����{�GT"��l���;_�M����=p��FeH"�6Vt!!Q�#/�ȵ�\�J�f�0�?Mvv���~TmN�㋿��ƅy�m�X
����3dx��Z�Nm�]�
���mY�p�U�[�8G���߅�>Zg��^9}K��{����ȩ�?�_fB�+6
���~|�S�q���'
+�P{6�#�@��f����T��jeg�T��@������l�!i������H�G�S��~(h^W���h���Jo���ZaU� �5�"���o�D=��r��-�ELN�����mMeY�ٺ�u��96��B�M�А�;�"�@_�������˔��@H$RyY݃v�"W2���(�˻�1#��W>e��u��Y�:%���"�a*�`[7�F�|@?��7dE��7�B�
�: z�7���u_A�I�����u Z�.��Cs�gP��f��J��(���!�淣I�/�{�c��J���D4�������g���e��l��^��o0x��U.t,g��,�>*���$�~�X��<����2�/��--�ޤQ�$��=��G350���$WÈ���#)Z�5�g�ݻ��J�"��p��:&����v��g	ӵ�@�d"�%���f2^��3�!���@<(�J�E��d���R�����Osɶ��$*2/���~[ �wJf'��E$1W�+zj�X�, Д��1����|��Ԫ��90?f�lg;��݋��N���d�&3C$F��Eʢ>�����kc0��޶�,%�E�fUD���p�ڶ�[��`������,Ѻ5+���-�i�����e8������ܹ�bq�7��hA[f�Z套�Y!/=x�.�5"L��R�CA�^�K�(�}�j� ���&Q������ ���$��{19��1����C��ˠ�^Q���(�j��w僽�H� }�/�}6y��8��/��wKie�;��㹆�W���'��b�Q�cJ��G��0��YM�L�D^r����_s�b�W\J��Q�����|Bsjg�q )od����&�ސ�+��P�by��
��&L�`#]�k�J���r=��	\qWz�7	��[6x�)ߦ���s����-n�e��:n%�;�?yi4և���,�rס67�zo4�Ё�ͱ�PA�5� �����������1�do�*cy��YgIÃ�-h�*����O �=]rDw\�n�&��|,���,C	�1>�T[l���$^/�oц�9x��M���׼n@��M�m�?�S5ԽI��)c�a�����B�%�l��6�'ѓ0@H\P#􁭏7X�ch1�����A�o�lX���	jʿ��%�*K-2(�� et#�Ϩ�j���������.��z覰6qC!
MZ���B�P)�Cյh�T�Rca�Wp�C�+*X�b�s�U�,ŀ�i!�/9�3Tª�����k-DT� �'�����-�ݢC�ѣ�5�,�~1��2k֚��rg*(ĂW��l�O8�혲�ɏ��p]���Ma|����l�,��U��N�r~��W��q���Q5H��ސ������C�x�[g/"&�_F��3}��y6��Ar���6%�	t0*z*aϟ���$�%��v'ƚ��N'/��Z0��"`˶#6`!s5�g>.�u��@@f����>�h����A�ކ�v/����i(��ʀH~0Xy�@��@:��(es̆ ��ɘ�v':X�S͖�DwO6��1A~����)��A">�8�Λ7��:�@Fqv���?h{��� �d���00&ۍ
2��+�J .���B����ڤ���cU<�����W�<������u�*�>U���ntr��Q��鬎jZ����2j���e�� �A>vf�z��2�ը���ߩ��"�:��?�m5�z��z�Ȕ>yZ���>g�:M.�׺Gy���'�/`#s�Яe�/>��U��h	?����9�P��� �q+F8�S��1�6f��!�������!a y8z�j�͈|���Nz�q��'\$���\S�bt-�[�>{u�����
��B^8��lA�!��g%��^3�5~��m��a�E-!��VPi����6�{m/☧Z�dLE�8#x�yc�<&���*���ܖ3$�X!��0��1��-��t�A<��P[��fr8f,�$��I+?�8���$r����Z�����!p�tx�Go�-vܦA�C�l�j�P1 y�C���?kכd�	�ˎD�A쨎	4<�������.x���b��n|e�i��M�V��uNt�8���a Wz�a���3, �H�ӡ]��?ˮ��/�)1�6��kۓlV�(+��Tb}k��ox�F�955,���g{�&ۆ �[�|\�����ֻyM&_���������MlI�=�����i�-�	�������r	.����A=^��򜴇!1`�h��~�2B��P�����M�����-
�ʌYO��@8i��GI�%Ƚ��A؍7I1��̇���>���?~��м�\��ڣT�kz,h�{��)͌�^cRH��t]׸��m*�J3b8�6d����-g�`�@ڜ#%V��*�s�=f��T��^)�	�m�{l��i��AcSQ�4�8���8t�뷔������LB�ο��y���}0�yX��Љ*�.}9�"ή��Lv��mV��q����ܨ߲���PɁ`�D��z0�[v�pc�oٟ+��$i_�ʉ+FЛ}NΧ̦�ؔg��>��v�'6��<��`��[�����tѰv�8��
��a�n�����:�܀0���9�(M3���i��d��\j!�@��(���/u1����:4�K�X�`���ff�x����P�O�w��h�-ڎp;_�7�1ɹ^�|`~�H2�������H���Km���R��Q'm)��08=�4�?D�3*0�2����W ��#?3����3>�2��j0_c��o��@��ث�7gJ&i�z��g`�c]Db/���k��J�rv�+ʟ����m����"!wQ#�M*̒��S�)��$@ɌN�f�%cj0�c�~�Fr��7f�/��P��DHJą]L����; �M]�"K�|��m����m�鲅Et:}9�����{FE�M����I�h����r����6k�^7�)�v,<�����ֈԽ� z��AŔ2�z/�z��U�#�uM)>��n��3F��g|��ְk�I��.�
�7��Ѿ��9Tߨ!��p��m���s_�(�9��h��{������!fU35	Q��60 n�����>�[��ˢ�Gb���QEqs�O�q�q�Hd3��j���)�5*rwn;�U��]{�Xjt���qAqu?B|"�ITx�`8���H������X-�n/�ʘ��'����tXo�H��ī��`;{���K�2({�蠙��,)�Ԕ�����1���d���B����h�I�Ҟ��dN��^�"In���������
�
%0�x8�a��% ��y���u���ӎ���=�0i���0���u�-��Q��2���$#��k�}�ڹ�;�����NB}(�r�-����k�
�*S�����$�h�S�*�j����B�:�s��M��-��qz���dDe-���S���׮r��u�=*_�!B]z_R�kx�>�(�6K�h&]{�������#=�����:�	�4��.:�<B�M����t��	����ѱ��ɻ��[9y�7#� �.\���-hD��[.����,�0�bi��&�/�i���,�p{�tx�X�D�!�5`�÷��g�aG'jP���:��s��7��"�Qi~ �袛��j��9fv��i?y��,��%qR��I��,V��ݯ[��}E7�����cj�!^���d\��h!����7���N�e�u+0W��A0��J��Ĳ����$_�M��]t�����+}WJ>>�5�!��!���2��j`U+f-��G���4�I��xE �e���!�i�k�f�c}p�=�w:��jE����%��z�L���$B�V�e��36��>P����~����s�d ��V�u���s�2�d� ����r�4Xʭqk�H�~��YFȒd�0)���v���ܖ�7�O˃�~]%�|�S��us����%�v_��s��� 3���	��1X� ���w��;�����4U��R���Ǡy�"��%��l#�<�g�r�z������S�1ߋ�5UM�Y
(�}���?�Z��B��dP�� �JB�DI� �P�P7�c�&G�T��5>�����Ȧi�;m�t�`�]����N���s�V��qˆ�?��1X��IL�3�OZ��E�p�(f"��=��韙T9�UI(ʀ>G�/���/2�g'�ѩ�?�%B�r������*$��.�u��=L�E'4VN�0a��$�e���	�?C���9��z���K`�]b��H]NC;3�F^�?�L&�sBsshΤ:b�c伙ٯ���=��n�l�$��������С%\�����4�D�H�G^d�d3�XF�M��&&����{� ��q1^d}�ꢹ<0�ϧ5���J�[H5��N�0&4��klX����@C�B;�;+O
���F2>D};d�Gj��C���yÔ���"��Ȇ�:�בּ����_Y�a��~������+N��Yn��ejx	'�Z>:��'b���`C8�=p�@�3�[r���o�(��O����Bj�Oq�b۸��pv�B�F�~��1��y.nu	�U��z�R���ꉻ�,�_|�4drc��;��c�$,������N�.raʖ��0��n�`�A�F�L�_d�A�Yŗ1?�R�ݻ���D��x@�?�9jqW�ʎ���'�`-�DTe�h�i�D[��j�Vsxx�lS�dS���
���5�=W_�%V7HP�^P��f�O�����X�p�����U�%�F��(����F�+���th������T�௘��]Y�7�1���E��ɶ���+���(Kʤ�%J�w~xO�iO�q o��P7��� �/�'��5e_B�R� ��� ��˭.��$I",s^�;ʓ�2I��$Ǽ&�>�/q�pn��m0�$����K5����xE�4jTF5*KN�5甖5�X��N	�^�#/��+����F��hl�Ê����c��fJ�[�G�����-vU�V�KI<���n�#Q�}�ˀ����f�@Tp�/Xz���k�)sXJ�9-=��c�-�):�:���6:qS|m4��*�r_j��䵸�18�ӥ3ZNp���R���+B
�����:�x��[&_|�ξ~��$���R��/!n ��L�"�2n Ǌ)��U��Xe���t-L��aJ�,��h��ls�߾Y�+���%����� ��ӽ�VFO�8sM6��6L{��^޲�������GA�lùK��	��Fž�(:!$�M��2����2z���%�C�\��7��;^�"du�<���:��ж�}����xǴ��\-$[j�Q�i��3���(��8ջ[���a0k��+�K�R+Є}��(�+Kb�h�-�� pۋ$vL�Ǌ��]��Eu���ud/_���O���c^v��o������r�Ϣ.xǛl"ϣ�N�:���Ӆ�u��ő�Z2;E���X�=l}1I
��4��B�Sҷ�'�9̔m&�\��N�S6ظϱoٯ�����y��M��uy��!���� O�"͚�bF�gG�aǮQE��%�K��N�����3ji�m�I#�̃�1�������M�Q�X1@��=Q0˯H�v��Ҏ	����KM=�}������@�g�1��j;<3~)��Q�Z���WQ�0��mβ��XW}ȍҮk��8�$��j��0תBL/5���d(�|XR���/j>�;nOi�G:�Pm�T�Cw�'���g9t�n�j��ڭ�������IdQ�S�d��(����4������U!!o�p�q�E	P5�����[JF6��r[{aP��
|�d�P�\r�Q�Ӣ������6';�z����6��Kw�P< }!:s�3�Od�?�b� �+�r�̻�nl9��毜�j`^e6�~GĜ@\�I�D���tiL���UH��&5����ך�����.����xpJ��iP_�Z�rL�Vπ,_���\Б�cؖ�$U�n6�v�J|S2߾�P�����%����AXO
Ih�>���B�GI9�1�s��)@�&�w-�䟷�y����ԗ�����`-r����_V�t�z���:ln9`:R8�'|'D{�]����j6��T��<쩉�Ҝ�D@�͗�Xo����rx|�rE�Kp��J�#>S.���"�$�n����0W(}Z��e��sN�`�I��o�x���
��ʞ+�m�J�*!��ߧĲ8�N'"&&�w4fV�Y;�
�#V��a�k~��3���xG_��b�}�N�;���� �U�5��k2���rl�;����+�5&���c��"(d� �0o,#� d�&.}�fEU]�LG<��O��]I��r\Y����vN.��0�t�Á�ۛ-;b!~� �����墭}6�H5'r�_X*��D�z�׀ش\NQq�.��^���� ����L]㋄�9�������ߎy�2����M[Аɖ���=��b��+�H�}"+�睝]Y0�1�f������5�I�9��oH�Bx�]Ǆ���@џ2��OO����gr��C�G�m��W�l4̮`�Ea�L�%~�N�ܭ�ɒsu�DV�c>	��ڙ�"�8��O��3ǧ$����'�z
[��ǰ}��]+�Xچ�^>��
JV5ٜ>�&@������)T��͉E����~��e��
�-7���Z��L��we�!��?��q^�F��]?�@�l����x�b������<���"�p�	��]]3&V�rpxw=�){sV|o�@ŧʊ�7��y:Z@��;G�� im�,%R�eT?Ls>srt<"`��s1���J�Q0��+���^�%���Nk�
� �����k����0�w��X,Ls���.O�(�z���u��WR�wb���=Uc�n�3��Oke������Q�5Z�g��.+��Z�����<�D���,L�'ݸ%C�������ZL�K��O ��f__��bl��t[���
���C='u)K	-W��Ř�6���."�	���[��[��<T(��Fd�^��Ȩ!��U��xD���#�1��#ċ�'���9}�8�ji��EvDe��	<,�:��X{��2e}�ĦpG�pmi��!.�!`C^P�`}�:-ڱ�"�rK7+�<�vb� ��mQʪ��q��?1��&O��k�MUWn�HS٪���G�`�Ѷ��|�N�v GI��EO�tكj��c�����yR`�M؎��g�����[�agζ7x�"5J����T��"gy�����&��l�S�7׀�����N�4���8q�`)[f`���]9�d�Ƿ�R�s3 x�|���}��/m�-��XH��dk�	ã 0#�����"��CV�I��܋��k�K��=M'�g��z�]�#�އ�o�8��u��\#x^�f$^�B�h���u� i�>�f��}Ћ*,�4ǔu%�u�d˻�O��W&����
s�	�y���i���;P��wk�����R��&��s�m�[Z{�h�Ň�;YT`��,$�Dn,���ix#�"�4�_I���uw��2@�^���b�����#�Q�����
8�6��gôe��Բ�Js�b!�D�4�L�-��]6��>��r¼��,�(N�k����$k���S �{M�]����?�����{�/����&�L5��$o��:�Ξ��4��>�/z�Y�'r��#qĥ/֦a瑎�eW�OR�_�m@l�L;nt)a��rb�Z#2�Q92W�����W?�����H�:�lWQ5w�X|�U��Qp��M VmS�5~�kZ2�D�`KCT z��=P�N����>���>]�N��肹��u��~n��f��hS,g5�ޥ�cZ<OJ�P��ݭxB�\r�O'��z4M�^��^7e���ZJ+O:��B��p]��)$ p����B����}s���QմK#�އ5ڋ��S��(S�I����mz�N��K0֮~�<7<>]"'�N�U����v���$(�{2[#�>21U��8Nv$' �6��_�k;4��p+Я�K:�����zb��G�`C� ֒�� �,�F��K<ke'J�aX��C¤C]���zt����m ��T��sz̽D�)�,�A�q+:���v���h2��v�A]m0A{u��5�#��r�zOY8:c�;:��/��h�4�y��O�:fF��6�O�B�]Q�̆��m��H��U)4�̢b��[5���$��߽�v8Y��t}�����B�my�wڏ'_�#�;C�B�WP����u�9O��O<t�.i�(D|��(���}ڍ^/���m���I�jt������~D��	�Ձ��y�����1�Yo�(�Pi[�$hD&ϖq_�`�Q�2��-��y�3w��<<��ڔ6Ͼ��ѽ%_	4^��FƂb�qK-�kt~�ZU�]Qs2����s��y��A� 7@���1�x�
t�	'�%�F` v��S#��W�V�.걛��jd;c#�6#��N��֒C,��	������""��[�驧[�K2�0��>�BC�x���l� W�b�Z:3�º\F�S����+�=&�c�/��qΜ����pR��Sf^E.o�4���7U�v�z�Lvıs�*A@_ͣ�K�ae9fɜ0�D0J�f�,u#h$&~��Θ�h��XK��I��̦m����M����
��:���-��#p<�������V�fѸ}�^a���s�CՎ��c2��M��?�?$v���wҌ�;��Gn;bGHނ��ɧc��j*i��g,��坝T�������I���Z�>ĦRo���z��$hg5�-�� ��M$�}�yJ��AH��C*~�ʗh�Ck�`L$�K�4j
���_,ϒ�8�F7��ïZï�kdz��7�H<pi�� ź9�_"��Z�Lk~��5E	�0/�56 `�~�!݋�k��[aJ4j��w�p"�T�b�'���]QĹC~����&~�k�d��
�QV4�j��� �N^��M5���lΓPrG��Q1�,�$�s]|�O�ߞ�����v@��?��7�����<�Q�`Cz8F��d������,�R,��J�1�� *�X��S���rh%�ƺ��s��M�)������=|�̆�������q<CS�L������5h�j��GސF��Ô�5���-�sՌ�5���g�s���bڒ��0j��`��� ��AOM��_Kkza��%'p����&,�R�~���#�p�E�hQ����Xz���Y �	���O��M �����4������MLu���סGa�XN��41l�ɥE24�r��}���6Y$EZ�H%PG�lX�{�qqD��3Z@ã3��}txvS�>��-��Tۇ��)��zj�w��	wu�}8+�bsƜ�O�%(�\[�'Kz�/� 8X�C�D�rڛa�G�\��Ps�;�\��@$r@�����=X��|7����i3�\ *I�s��k;�G�,L~И�����]rP��..t��_�z�u{�4�1�����vF�]�
��4i5X�f[ǁ6��P�Q���Tsl�U})+�VjI��|ղ:�W�+�҃gwzo��eT�x6���X�v�mZ�4���T�����a �D��չͤ3=^S*��x �3���/"��Mҭ/s��&KG�r�K	#a�}�:�|��/ã��qǹ�;/�3�G'�������MZEɒ��j#95�LR/0G��9��@�Yr�c��l�0`Y��n�,7RY��\9 �4stH�_?�M�8���vC~f�࡛~��C�!���˺}��.#�ɷ�!�����d�[��S���v����;��3�d/P����Q�J�#��!j��ǻ��FP�}މ��ĺf<���A���Z&�F �����-HX�qSng{+15鱍��a��׮P�"��o�ŵ�����i���c+��R����o6�m_M�� q��I0��^R�U�3/�E��A��Dz��¹���,�l�>���w���0U�<�"3�U�5��?v'�@�wt�<���Qږ��'�1������/M�E�a4'fP���r�?z*�Y�
�9�-������!8~��4l}T�K�ރ�e��?�h@������u��ļ�x��\jKb���R����c�^v���ْ�Պ,s�Q�T�xZHjQr������ۼw�V6�
������q����3ﳿ�˩
�7֚��=e�<����=�)��g��^�S?��n`�,d8��\jS�Hy�h����T/\�/����
#�j%̱�p�������+�Ï�z�N�^��N[O8�p�,�h�������-��j���y��]�9��R�R'������׎#���y�X�)��v�`���TeW�ܠA*Ӯ?u	;W����������;��_�i������&X8�/��O�ǐ��),m,'�(�s�.�Qk,�1�.$!��S�f�th�QM���q���7��9g�-'�9�����A����|�bt�E�Ua�W�^@C9��B{baO��WJR�7$ܐc�C��j�V�A=:�|��gA�<f
�B?bH���1�`��nG�{ED
R�ݠlN��rx��p��r�?(�Qt�������~���$Zx��p{׭�dĩ���VǱQtݚ�&�-e�6�����"{W4�?�]��Wfp�L�5�疫/�
Fg�{3Z`���Oy݈��n�xy����k�.��h|�Φ'-�U��K�1�z�u��y�e�}39R�&Ŧ�� ��&�W���p��瞛�� ����O��7s}�	-�g��}A@|���M�4Xߞ�2I��l����12ss�G.���LL��}�/������L�97��?�,I)��$*� ����ƛ���ɺ�t��=��C�B�9(K�u�jN%��*��L���I#��Cv�x��~���`ZYף��'˩�����Z���>Z�U��x�K2\�U��7�/(�~�q��aԸ	-4����#�l���PNiD�If���Y��k��y������(��-�8�����'�^�����bX���p.�:��E2�Q�f�7:b�e� mi��^���,n��q��pD:����4y�i�#�3�rS�b��{�庴������Y�*�9�M�m]^Twtr{����qa
���k��īev^��<��D/9�����:��T{H���]�E��#Ew�m����]1�|�c0�����G��ļ΀ݚ�&*�6�	[�욱�-�CP���ɉz�F���o�b���<c}��X�4���a���C�Mێ�D�L��h�L������P\hjY��4�bo���a�b_iw�Ju;*��Յ���N��ם�ԕվ�@�2��
�u����,����͖��#E�`�&Ќ6�<P3[#G�l�l�6�������#E���^���vF�y���������i��y�r^P�ØE�!�����x��b���װ٥�I��$#��V����N��2v|ae�Ł�(��22�Ə��aL:�I\�u��!�_�N��Cb�Ϛ���k�����7'�V����~����U���07���e-�'�j�W�M �0V�ߓ �����ظ�0�����,�j��=!)����z�6�.�Vpb>��J#�D�՞ɼ��&\��O+���:˅ 1E����_&}&�4�n9��7���X�Lj1A�O&��o�b:�^�*[��p�^K[+�BPA�d�i�\Lb����=i*:�WLb�����!�H�5��XчGcc5��l�(s{��J��d�@)�:�{�/rQ��݀o�6�r$7p�̾�˒����"r�F*��my�0AD��B�V+M# ���X�[ۿ��T�`X���a#��?�m�35�e���JS���Xj�J>���Қ�WMD��;��.H����l_Z�@8v40����C�BM�5�sD��X6%p�gC=�w��#��ԃZ:{Ң�#J�+��L(C|�c��d++��>ݝ�����l#��SA>R"�7�9֣ç1y�É������3�<���#�ɐ����?���D[���:����.���N�=�!M����묊��V�sf6$�͠[��Gj�}��$����s$5�B�NTT~;QC�������Oх<`SP�_�ξ���&�����K�=�bA�Pb<���C�đ~#�o;����1%����nj?��^�b��A��/��`N*�*ː_�Ss�@�KQ�+�7mM\�����mF��	E���yE��F�E�?�`}`�\G�;B`�8�07����`R��P>�����x�����cH�8;�ǟ�BZ��&��L!DH�K�N)��L�C�� c��,���dv7X�Q�&�\�x���±ʹ��2φ+��	m�D8�~VW��9wd��s;{����j=�Og���k^��v�Jͥ���1TxLL�r��)�A�F��k��(��d��OT²��^O���8�j�35����~͙�{K̟?���x*mi���F�����n����ܬZ�,⊒���g��*�~�`r���Ý�$��s��b���ڐ:�8Ƀ��sE������Y�L���3��klWxB�y�2?'�iԻd�Z�xcn(�'9���y������N�W����?.������Uw}֖C���7��m���b�R��S�za��3����@��v 3pD��8�!"���7l
���Q]��ۡ��*SnCuR�V�Ò�`�����˶M�w7-ӆ����ԙ���ﰋ8j<�kPU%�1~�L1��H�����r�V����&9�s@ɰ[$��xߥN���lc�EO^����7�Sת�Sx���g	��,�*��«��I�v �p�\�J=ϐ
#s��@���f+-b$�-^(�&��i�z��S�4^�,��䧞ȳ˝֞� Q����x���5*��#�4��Q�J^W�K�z�7`\4�x'���Mn���"��~�8W!��%kH���y}������1�mE�,a-��`w��*�nIy��(���Kv\!�!2�� ��mnR#�"��]`:�����D�����fpaN�'�2R!$�q`����ʈ�ѓ�k"��7�W>����*ɞR�����,�n��x䲝����Ĉ�u������z�w�}`s}�"ؕ8�l�+����a�q&R{^��ț��@�壒�?0,���E����>����WLO�WI���(��������"0���1{�V���R�eJx���UZr4+���x��a����"=�#$�䈭��Uf� ldL[���s� �=b����S��#�1���Jp����r�/E��&m�ץP���{pJÁi�&��M���nc�[ �˟��C,����!��\I;~��9���@D��y'ĭe�\T	r�p����Z�f7�.���Moq�C'�����Ո�E$�P����ea����Es,�>0��`D���ύx�9q���c����;(l�by~�}:ZW6o�Yl��oXKFf�
ch`�\�j깹eH/`JKۗ��^����n1R�qY���6VhfbOZŊ�4�*�g����
��E�n��L�_(��c���R�|@�3�)R�_��@�4iF�kl�)~�ԏ�kT!t��|�b��"g/0�74p�E=�^k����{XkY1���>�NK���2ARv�n$<��	"�[��ڬ�5�f��!��"�	B䚔��������b��>�#	'!�����#��zw�~P3�0�t���/����B%8#��3�C����`͈�.�N^_SUm�����r�5s�c�������`rl�,{�3]��#�O��a�S-�F�	�<e&�0p���_�O����Z^4|�ޯ�y�g�0��^��vṆ�{;�CBW����l��y��D���·_���+�U��'�����PA1�j�nz�_/ÿv��G�i#ߏ?�c8�Ę� �	��l)d� r'(^��e�8?f8����.��Ԅ�LKr+�C��'7g�;���v1ģ8hq�Z�m��?����:��o��H볖��/���P���+�4�:�[E�O^��g�Y�9���uS��������0�'"�־|���NA&S�<�.!��=ٛn�D�.j(�r�9�u7պ
�p\k�ؔ����o���O�o�7}g���0C㫧|�Q��b�G/�����8�����hAV��$�t�_4�_����$y�Ǣ��5��ժ�+9~�>��G��a�$� A���|��!jJ������k�%�Y�r.t�n���<����:����B<��QS]K#�m*��b�����\���&����?�P�/�{�Sz���y6MM�K ��eg��V�����8��M��EnR�5���{G� �}��H3�N���7��Bs
��Z��aH����~�\~��脵�nĮˈ�HVchN����-�K���l�� ��A�S_n���I������e�w�	B$�x�S��N	$��|
��䑼�׍��}���(~K8<.PX�����A���Ҙe������
ںW�tOfm��j�r尹Z �����V4�O�b&�������0V�J�������tQf��S߇�A�s^
E0Tƿۣ,fI�x�ϔ�cЕ��x�����V�P95fUp=�=��w�H"��u���A*��-OO���ރ���A����P���j���I�S~��ڈ��vZ=�Ue�`˪M���d�Zm=�\D2bh� W:�X�p�0�8%v�E7]Z�1s��K9�dѣM(f���<�t���B��Qw��+����JP+�_u<\n��2����:t�M�*-IC�S �����i]Ϩ=_q����'��/��ws/����,��b��Ŵ�Fs��'@��bM��x��ϟO��B0�Dk�eD 2�ͭ�_��	�vJ\y�����<64�*�͏<܊����	w�L��zseWD�LB)�6%��x(d5��H����N[W���̣�uOL1���������4+#�x���L5-�~k��p��ZZ�[�YsN�+d����!RS��%:Pa�1�M���OMG����w	���0�a�HE-xpȾ�c7��w{���Q�X<����ˮ���]�&��!'��ٜ;�����Q>����p��pcy�u�L)����r����E������)ŐJx�bc`�7K�΢�k���^����w��IG���m��¼��Ś�`���(b �������+0Th�
��5ޖ�Dk�Z�R���F/
��H)�W:ۏA�cM�km��Ny;n���c���a���m�Uh�����93և��LA��QL���(�D`t���2�{��Np�Q�'פ�R�ڧ1eYg�+��$��TG?�V6!�m�����ZV��7	�М>W[a��'�!w�?���hŲ��ؑ� b��0�ɦ������ ���$�����9"��ꉬ�d� �Z�9�X��셾?�̋�N��sP�jzl�hjE����N\�ݧ\�c7���i s80�'Q�Z���>��h���R�o���J��U��{5_&���Wu�\�"�<iǍ��ϰlg��'��O7��6r��l'E��Vgp�������R��H!�B�	��������53�tFCU �[��$ǕH�;`k�ު���=ј��_����Ќ�SX�3���8�x������G����\�9��$vA�';�/�5�Q2��=���1>�.E��$u�zw�C� �IY��R��<����!	�G���{�?��~���*�մ_����w��v7`��l������6�U��c�+�<<�o��D�	x��IN$�p���� ]k���M�
�k�pt��?v���`�߸1gݕY#?�8�0�B)��i�q/���l�ը�/�#��Yk�������x�)��ظ]M���	2B�+v`� ��0��!{�6���!�}�����
ۘ�f�0��h6io^�"}�(���8Q��\k0�`��o`�?��<Xm"��%�f��e_��=&^?��*�3%�fg��?�dvėζ�%�n��i݁p�T>";85�v�"�m������ԋ�^.[P+:J�$�<�C}�:ĥ�?CK�Yb:���a2<M
�>�\����
1[�����t���R���˩j�[&�ƭ�4�^�4���� N����
ҁ�ꚠ����al-�ѝG�f�Z�"�ݐǢ���sK҃0Ur(��ݰ�0��%jk�ԫ�1{�]�7u"�8G�Y�B���4+bm��p��lؑ�N˅�\N'ғf��I\´j ����A&�"u��[�+�}��υu2+$��wG�'�
Q-J�m�����~���sj b1�pحTqK�� <��.�9�5Q�;h�&i�Bc���A�g�k�f�UZn�E��K���Q�A
�2:���g�j�g�7����I��G�$k�!UJNU��/��[������u�#gJ�7+��)Y+X��l{�j�P`~nq�8��⧪���v�����	���<�j),gQ;�
�I𓙋�f?����ٿ&y8䂵�v/ bmfR������z3X���#���vl��i��y��
��Z�7�V:�� �K���(T9��g �5^����)�J���L��$�d�f��J���`;�8�4]��P�#좶���!�����)k'��K �rظ}��8�2�o;�X⡑��������`
�vc�}�
d3�k-��a�ev��;��g��N'8~D���q�h=h����Q�*3�W��T_�s��c��^N�xމ{�j����{�P>ղ��y>8�{lr&Iܹq��e��������U�z����7�.*���l.ê
������ʬ�F�;�{0�1!�EAG 2���N�(����p`��η}���|��.j%���{��9���p�(�[���
Ady�}p�+� Mz�+i���{�b\|�c���1*��V�8}�]q2R[�*���&�  �TR��'�+[�~	#+cW�~0N�!b�ٷu��/�/@�=��5�lr�MГ�՗���6�V��u��D�^5���I�M����ށ��:$�g��K�{�����E���ec��BC�K�[���6�Y��nB��!�E�J�p�[�Y>�Aw|���G�8���/�x�&���m�����=d�½�A�ij���:�I��(�PD!~��dF���i>W�m齡�o�˹�x7	�V� 4��؇�Q�C 6<��nQ����� ��]�Ѹ�=}����. 8���I?�Hx��:��k���i�{�~�<-���d���'8�>K�50W���ɿ������Ċ��mH���0pR�++I�]7�NB ���s5�qҒc���N��3�O�&/��%�n�V:�!Z�s�]^����F�j���'H�@=%������L�|/���د[;lf�Q�v#����g�̝��9���2Pǘo�"�q~)�:�ٰX����EP�����E2m�T��f8I��6�>F-CC�G^�ֻ󻹧�cp�]H��������l�ywT�l^�V��z�I�Y�κ5f��W��:�����B��?D�l_Ӕ�Ӕ0���Z=�$bu��ԋ5��f�Os�.#FQ��h��67O��,M�P�Ջ�ZY��:�L��������2`h�w�׸7~FR����"^�G�v	�\�H�;p�c���U�rM6G 8��y�ޣ�=�/�[�!<���YIPJ�*4J8�h.A�XߟQ.w7�[^L�)
"y��r�v�/�ͪ[��$�Gs�!_�Gx� #?E#��[�0�5[���pW	�-N��q
{�$Q"%s�"���T���mk����F��e��f�p-y-������Ϲ٦�Z�iN��"��D5�f
~�Mh�� i�Cm���@���xdi\�D~7~�l
���s{hv�Kn�����$��SE"�����:�ζ	T��p<�EN���({ ��Lx�	e��� yɣS</��>��N����8kUEs*X�j���[A��^�5c��"�$}W;㓩#�_���Km�~�ˌ�����5js����SN!�����dz�#��c"��iͤW3����H»��E���hpò��؍@2�/:(�Z��	�^�i�#
c�ֻU�
OZ#ޕ߂�䛺��ʧ9��w¾�I�,re�����\�����י�|Φ9�xC�>�j����N��SD�FJ^����]�ؖ�������4�����B�^��]\�Kg 4)J�Z}l�"׻�j�bG�U��__�l�Յ���%�Ҵ��<�u�R2�v�O�e�<Ӓm-�&U�c��?���Z�&b�=�ה���!�����~�"��Ck��z�C c�R
��7�^>Z]����� �]~��+�4 ��F��R���-<$!q�G4c��(a5Z`!�����YC�XX�'K��t�(s����"}G��{��1�_D�mX:��>,;ѱ<�����|�R@UH���e���У��K.���ۑ�t(��z�ֿW/YiLq���B+�Ԫ>z��vC�;.��b���z��L�F.{ÞԈ��m$}�=%�|��QU]~��6u��c�2���ڀj��-#[�ΩHe0*k9��g}z�}�%���&�{�梸8y�H��A� ���!٬֋��AF���ڂ7�CL��~II>�ܬ�/�*����k��� k��e�W�\zGS�&Ṙψ}��mj��ps�@��6�(��Wdd=S�X7tUy0�n��SE�H%_�t���)�Ds�N�*Y�?����6 {��`��=ǖ�W�����m��L�������E���5x8�i_m#���>�E�̿����|A;��裿-d�u"-�in���������_q���m@M·���%�E���D��~�u��:Ex���ܾF3�#��9�	��ܳ����-Lt�&�'_LD^�]����H��;D��m�S�����ca2��>n!�1��w��=�aQ��m�
�~ku�F�bZWI_6h�	��P-4Q?�"�u��	Ů:������Wv��]���\�*�ږ�0f�~:7C��M�$��jH� ���M�\�]~D;t�z�k�8gf%B�Y6�~"�C�x7�?����a����08[�3՞B;
 �P��reJ�d��?!߯!Oࢸ$wʅ�S#GGE�n*I�l��)��*p�}q��
8{�t
x&~�ZG��������7��5��OkY0t ��:X�3�ԍYb�i�	��y�T��G���5pn7MMl��s���o��̅��$�
�E9�p�i;E�Ulgb8p��pڼVV��}�x[OF���6˞�q�኶��,� �T?3;N�o ���j`&ǰ�P�Ɖ��}X��MF�y�1L��V�̈�V�꼨�''aW a�D�io�� �͍�7��Ye�x�Dk�s���$j&ab1L�V�B]-�"g��v?6���V'~Q��^j߷��	#�wא��!:BlZ�9@|��vd�#
�@v���C/B�|-L�� �{Ϳ ��~�7	��0��ox�A�m��庅9��ެb�� 
X�����$�]qg�:@�`*�g>�w� V9��h�qt$�UjDl��$F���Ji'(-ޟD����Y�|�9LSWQ�#Dm�^S#��C
�a��~^�h����8rC�q�����xivf��M�JC
Y�/#p.�y����/BF�4�C�8���"���e�X�*Ο"G+�;�� ����aր��M<E�J#@���w���傇���D��	K�r,�K�~�%�����f�p&`�w�m]*�Ϫ���Z��K2Ć­tM��(��q�+�l��/�N%�0��#�[�&���!���U{���|�m��E�Xl|��8���y�xIb���S��fd8����W��ݝʾk��\��\��~�9�yj�v (U5�]Q�9��f:a�i��y�Ǡ�oĐQ̘/f`��9��Ԗ��.X"1�������@:�"��/^�����g��'�2V ��HK���V��w�v��uZ�#?�%��X�y�
�*����8$��C&�B�c���	X��t�+ISί(��H�on�UP��jtD:�ϟ�k �¡��h�f5�+���NO�X��zGez��=��כ/Ц���;w�H�B#�B��O�� �ψ�!YeIh�&)m1��"��� �Ym;W���NA�	��.� g).���<�{ju	�婠�C��v{8�g�%o^��k�l�n��Q71S�/P�6�DT'T��R͠�a'E"v�������������Kn����@��f�B»̐�n����MK��K�羹W%�U�w�З��e�Z��.&�,z�Hc�U{|YZwŌ�9Ai�� n��馊Q��'[�܂�I[�IJS��ҧ��~fŤ��
��6��<�B�3dqIv�����Sj��U�1���C��%��Ԓ���b׺�.}�.��ޅ֊ݮ�uZF��e�b��+�?`��,'#2F3��5iG{��^��П"�����X�]WY�5�m-gBw��n���{�WSu>���V!�
�l}D�Sٚs�kl ������Ϝ�[���ݙ��R�ds��{��dt��V1���^������ZV rĭ�q$xڢ�7��v�}�eX�����!e�A5�-⯻*�`�24xF��3ۮ� C[�|L�?8��3�ȗ+ΜE���3r���[�Q ϼ�L��N0]�ühb���ײ{'z �6^o�Nd��Z�4aԋ9�s�^Um�� �xt;��Yx����� Im�hc�Ϡ�"�e�;yo
	ļ>\n\c˭���K�L:L�W �Shdy�_"_y*��`9/�i�>�������BO�!�G8%���K�3Q<�4wq��Ԅ�Ю���7���,�<mƯL|����12]����e<�v�Cj���@d����ǜ�
\<��D�$�$X�Ϝ� xk����§N]�1;�_��]�����>�B��U�s����A/�yJ�n,r�E��*,�~��t� <���GwY����@�SƷ�ڈ��EB���B��'�?kkϖF�Y�`+7�E��wQ�Si���W>{�w�<J���_�NP�f����&�cC0\�Su��2���l�/ ��2My0�ɪ�ɩ �A��3���dO����2�[=�/k�2�������v+��3iW|�+X{z]�_y�EYz��I�T��Ԫ��/�C89-�Oi��CcQ�|ĕc�/�Y����
��`�=���#+��]���E��.�]?A�3Ń��_,_�*�tW��y�k<�p2�lb�@nZ�U}MT����>��Άe��{�<�bІ�p\P[�N85=x���߉fƋ?D���v���E�GO4^ītz�����:qПD*��<o��(��7� z5�6=`�0��F�{d�]���d�LCe�:����Գgnu�r�n�*�ڕx�D.��~�|m�28�Y	���*�oN�������g�1q��t��#u8��}�%MP��}�k��S���WP}��!��'$�|�Q�H�ڝ�km�S�wlv�9�p `ŝ`K�.�K�* dU�J�
�"±������� &E����C�G�ˍd[w�����};��=c�OW.�[˞$���!$c��V	2"�#���8U݌���j�z6�:@�@ �|~�|��]�0cdf,�/�+�<ղd;���6�n����c��̿g��ޑ�o�+�B�c����F��W~BU����o�5t�F_؃�Md��R�c��]'��VO�OJ���7/E�����;aݎ7����᫁>,nFꃤ���G��Э2����	���^��Cs=����^,~	T���"&��YZ��/�v�/�6�s�Bbx�u���.ͷzܒ=AI�҂�Ԡ�Wk@���`�+=� 2�vH���DC���h+��3���*q�S��zi�\ٓ��-�'��M����[�5����w$G0%G�4=����R� *��X�B+���KN,j���U��9.F��* p�v����I�k^��q��BQv-���jgj�t��3W��6�53�����peO"�-Zo8�ʹ�+��=Y�8���T
���ܩ�l��NϳF�Sr=�Z�~Ц��XV�CuL�L�e�W7�t��Vv��?xr�GP��$�yȑ���% ���a�1���PM�u4���e�8?ĵ@�F?�y5�D;p��0�����(��v�b�����}Վ�:��2d�п�:����],F-gI�9��Y�}AF�V��#L�X�d�:I�l{����_�*y�c�)hY+Z�wF� $��'I������x��qTx������t�^������&*\�i| �"�'G��jL�&{�x�|��]�,�+��)Ke�P�.��L}=/�r����a�Ҙ�vF�?=�j�t�ใg��JO���5YJQ?_;}�1;!x�K�#��IM����jڞa߷�nV�7y�7��~��J���: +���N�4
���E](cC���Bs饜5�jOd��n����$�W�N�]���[�b���X������':�<QȫB ޿ʂ�k4J�Y^�5u�֥�@�v�lz}�{S_�`��?,&��r
a����1��Ot
$��mKw�Jnي��ŀO�����P/�β�_�����	�X�m�Yf�;%���f����DS�>�i��$����=���Z�h��p
�ٍ�S�p�W<m!R���EtR �ժp%���<��xv�Lv����b���	���o�����Dl�m9j�]�Z���k����k�^�m�\"���%���kG�?������4b	�ݎR�M�����N^lz9�˥� ��r�C�n~�ޣ��ƞN8��&�ѝ͈��B�NX`Ռ*������,�\w�KW���h�-kp�<��c�jW'Q��+�c�Qf+����]m[��
�g'<�أ?{L���i�˹4
��c����+ϩ՟@�� ��x�P�ϔ|V�:%�W\@M�
��Y@K:����?����B2B��de �*��L��uk4iX�^�H�nE��2u�yH�*&#J�++��\��j2"��`8����PG���t�}'��c.Q=��QH,#C�`Y���%�i���Tx�{~U;!LW��X�[~u��k�<�C�L�
���s�C���������NV�,�(jv�Z��K^~��F q�)R�,��z���:"�����ax��%cu��Bv�)��W�L#�{y)��nj�փs�f���'e$S���xdjhZ�<x�.�q��Mx��}N��g�c
���d3�Fr?�X
fC?������tk� ����RWC{��v����V��f�$_�X���"�@'?:��qN�Ж���Q>glɁ���Ykȅ����O���?~TY�{�t2m�,c���t�HM������#W�˘M_�ɝJA*��u��%9_f���63q����w����t�76��b�A{�}��'���@TR�'Fo���_�g��?Xc�Bw�\w�]�ZcD]���wy�/!�BN�7�9^�뗖'k�$����]�����v��^
�H�G������הq��m���u�!3�;��{u��NX#��8(%GR��E�Z���n�pՅ4�R;�����ގ�ý�a�ۇ[+��3{�������p  �m��X}Y�Ἑ������:���vO�M����Es�����L�h�E^�J?�5맄2ؼP+a�x���a��	hCy���<���i���c)v拥��J��p�8H�0c'�M�+�^D�8���Yk�z���7��؇�v�5�|�@���X]��_)(�۰}_t�p�����xB[�Lt�s��e!��x0�J�82Щ��*��������M@I�3�DHxysנ�-��׿�8{������ŎTw�6�c�u�\֯\�TsQi;��n�iq�	4T�l�b�E���2��{�BlF@i��������a\�]����Cu{��ґ</�>lP��f�L#�Q�7����؟<a�L�R;��l���^�ߑ������t���5$W�b� .XS���U�2C=1n��^���_���}w�r��Dq�'�f�3�#�S0xԂK�Ze�`��ol1T
a X%jG����L�;�d�g4��{~3��������f�?�Z6�m���#U$Y1p�	"QX�irB^�b;��۹�ڟ=a9"/׋�8���B	k�~`�x������O~ڦ���އ��PVlp��[B�r��9�xTB�J~������l���"\S���uO����&��m1�>� /P���W�θc6(<��|��uPUz�]�|ne ��V��h��lm�4�L9d 3�2h��ŀa,��t���(S��F����ށ�� ��o�w����E�ܕ���вPo6Jd&#�]}���qORK��O�
�YO;;^��ea|���
�"ƶD��5N�'�sFm��؀
i\p�רm���!Ԃ��Ks`j�0GY�}V��Z�#�(���%a�ä;�Zc�jW
�p�8Gjt	�����u'�d�މW��gt��0�%�$5��	U�IN:>#���Y�T���y�\]z�O��(�x�V:f3���X��p_J>R��Z >���%��&χS����*����v�D,�,�5:*'p͠ıى��wLм�?����`�:��ⵑ?	���i��ff�$���ɢ\R$��_��~��:�ִ���� ��d��� �gv�}8�����AQ���ѥ����H��᫞��(�ćVN�dߓhs�<w +���Y���r9�ے^u���?��NK�������c�g��Eyk��#`��PNnE��I�gR�Yv��`�t���
�J�  �I���**�G�1jQw��h���ܾG�c��=@U.ߍ�H�������,T�A;��C|E�@0��t��I�	0�n�2�sbQ�ת�%�b*����aIe#�dh!�Y�!_W�h �c�l)X�c̴+�M^�t6Ǻ|��և휂m�����n�Ϸ�y�`�ǚ,�4�KG��^5\���s�$D�u���ح����+�BLF3A�?����ۓO�����*��0鲾��4m�"�?��FH;ֈKd �G��*\���EaW%fm~/��|�@${�\T��}��y�Q�ˌi^_8�E�4�U��Oq�q�N��u���C����c��C��\Cxد''IvBga�?Z��;-X0�z���a�����u�����'���h#�c�j�[��϶��xd�Z�\�M'�ݶ~Z"��>���l����$�m��yZ'��{FEkh�o�kJ�!!��M���l44x�GЂ����������:����rv�'�B Y�f��f��^>�е���c��i�@��}if�ϑ <ۑ}ZqO�G� �6�x���T%<��CT*,��vz��#Y��UX��O�Gj�A�X�:�<o2�[�}!ε���1_�g���r��_��X�n��䠠,�F����4PP�j4uy9`V}
�z|۠3�nf���Z`�
�yHL�n*����Z-��.Dme."�>��������yY�?�)�a���	i#�$����W�/Yz�5�"p�҅W,�A�� �.�	a��$t�c	:������Z�:����m��M3x"�f��d�Ρ����0����|v1O��&��;����SS�M�w����������C�C��y���i<�葺�띆A�!���}.�:4�#3��w�B��!%��1��ȅ��E���|ZBt��E���n*!ې�;���lja���z�JP���Q�����R�*=#Bٙ{�i5U����.;E�ПT�Q�|�Tb�P3k�~������ȥeSiO(��rC_oq%�����s��kd:�Ơ��W�tt-���s�s�41kއ��Rd��?�7}�n����I奟i2-Tۮ#�����%)G&��z�kԀ�YƏ��A:C8�Lu/���d^���q����LiX��$z��꿮�XuH4v�;GN�+ʲ+Ŷ+r�#��V��M�V� �ӈ��#3���kmi�0���.���Ǫ<p@����D%�mp�@��m:�5����F>&t�����
��Mͅ�f>�.a.�.�]�:���	����a� !�Įxd�x$�R3�z���J�9f+�n��;��&g_#uLZ�IC����}����<<H��@����]ӎ+m�����(���bR�;?bb
��;E�k�u��7&�/<-r}� �a���8�uhW������Fb�s��7x�lQ9��9�+PV�A(�2n~�M�Om�A _��#��v��&�����/J�]=��Z<	ո����n�P���
���Mh���&���	{Dޠ��r;�� ���#�QfL;Ӓ�'��v�WD�Y+��
��>��n�
�	�O��?ܜ�#�� 	���n"ޝ����(�B5��l��j��k}�t��Lf�_+ �~����;[I��K7�'[J����Ŀ���v��!}�]w�x}��(�f!x��;G�Ӫ��-��:W��mN ���8��j����K���u�o�#��/���q_Qh�3N1� O��h{��
�A>�ie#8����e�r�.1� �|<}��vX����iz,=+$\G�̷���!���I�S����t"���J3��;D��^��l�y�4 A0���:�Ң�O$ƌE�yA��:��%9"�`�ሷ:@K,�ߺ�6�,LIHJ���y}Q��x'0��=����yHW�QS`L��?
����_Y�}�A�-~����Mp�O��SW�R���B[���x��q�0)�����ʯ4d*�p��������.�ə�CS��D'�����I�B Z~ݒ�4ҟQ������l����ԷC)u�k�N��a)㪌��)	X%��T���ڄP[k"�T�/�@�\�xpΑyq[y9�l��a��\���l��'0�E�?q*���3�o&��
	���	,F#���f߼m�qж�y�w\��Gi|£����� ����\\p
�����ts�4,Pǚ�w��dg���hI��� j�R�ɱ�Y�I�7�7�۾�&B6_�E�s�m UtA�i�=�	��cd�'�b�_3U���*���Z��1.(؍�^}�j���"4 ٚ�YA�aG��ɩ��� )�v�.1$���U�!P�	�ʺ��9���/�S��DO��Iu�xY�ԝw��P�,��T�,�a�t8<�_�w�t�46�IgO$��8��i�.U��ȕw�T�� �LOeJ���i��>�G�, ��[
5��i|��v �N����r�=�06�͉4P�1�+8�9���Cu��Ӊ����j�� �2�c�������v���.����W��b��j�_�b�K]s� z,�F�;�� �|�a����W����@����Ȓ-Me|t�R��Y)�H�x��⼦U�wR�vύ4����.��F�|��!�ʌ��@���9?�#���?���:z�<�of��dGgS�3NHҖ��Hxw�7_��0�[e�Q�4��� ;
t��?+�M��F�l��E{j'VTl����u��-�v�"ʡ��-
vf��2�q���
oh>���vu��_�Pu?���-����d�h�9�`�H����y��'��=���#ޟ7�%�)�k$�|O�
=��n��F�
Q�J�|�Ϧ,�s��&��+oO�a�k��CO��j0��B�9��[���B-��5c�q:?j�Ťz
t�Rn@��1Z��� ��4[��=jh~�c���ҖW�d*q�;����=˽���hR�<��#���'��l���1Y{!�&�;?�w�շ+��)��Y �]�scU("���;n�Z\��e� }����4!�����W�J��qLF'�[6�}�讏j�eC晨�C�y��zƍ��1(�{�2,�R>�����%�]�I�,�U�m(㔉Z���M�/jKkf�\����M�t}`���x������l�ʙ����:��8ݮ�kAۤ .�~�p}�rsi�&�.��^o�� �!���(�I{D�f����x`������{����6X��P
����J�[�3��)�������$�5E�F�x-�),JJ�KW���֏
VA�D�ű0�-6X�2^�/�]�pe�Ɂ��4&,���H�u.����S���BX��f>����q�����W�X�;e��A[N��,�8݊J����������q���̂��<�6a;M�?"�i�rz��B�e���/�C?�I��H>�nt���>/�Bcj��e�-W�CJM�45��O繆0q�e����
��J⯅�;|�!����#�Ǒ�aBz ���.���e��w4(�_ñ��p���$(2�7e�[����l�^��0
����Q�Ee���1̅��C(�Sg��S>�.|7t6��U�{^��2Z�
�G������4y�(����/sk@���r���a�>�+��PWW�|\a��I;�(I����g��3�z]���R�P3*C0�h]<f��h�N%{BنW�>�G�|L���n;�ҨS�⨖Č����=.^X�OFރfB�D��3#���a����-�JR���9��	�EJ�(�{ڎR�_�S��QןKL�xx	<�VƤ���H�:�yR,[�T�0c7H.�#b������Ķ����8Ǘ*�͉%)��eI��A$Rm`�c�����I�af��7x�|�L�4_=��!_��xݱA��;�qCø�(�x=_�q�}_��_�	Ǜ>u~��|���.��8~�ә	
u6s����A+L6���k��)�m�rqz��ʯ)VFD-��H^�E��KG���Z��gw��v"ڔ���M�R?~+
j�� ����7�-�m[%}���Y�����X}T�Q���\*�2��}����Ͼ��j7b&Ck�"Yo��3	�!
ln~�b&���nr2�98���o3!1�[��� i�s;s�ҍL��U�D��V�Η���N6��?�Y?ەJ
g���9������^�w�D�ڐw�c*S��B18v���ɮ?0y��.�Ϳ����ҎRR���:���j+q��̍���\�x�/$��2#d��3�쳍J��Œ%Q�!S�lv�znK��vm5�;�J�7ȃ�Ze�����	���{�.��6�,_g����"+	4�A���?����֡��(똤�e�	����Tw��| ��t� .����8����f5�d�N:dB"�_8!���}h���ys�>��K�v؞�
�G�v|�m���/luk��������h� H.:A�Ԭ�[��,��4`��\0H,�g��mO;�<�������7����k�4^k?ǉ'�Ul���"2]��¾֯�V�X�ԟφ\�~\3�U6�����ͧ��905=�>����8:��W���b4�l%���إc�P���R�M�u�h|j����ʴn>]����o}n��p9�$��5)�/Z�y}M����Rش�Hjz�"���Gz ޙ��DiL|�`�O�"�g�LN��e�4��̄*���?ᐐy�i��0�s�-a����=��Θ|��Y�+ΖJ�q��ALZ�c��a��F��
oѶ�M`u�� �f8LQ�+Բ�L�߿>�i�E?��n7$�$��g��d�۹���	��)L�"��xB�Rؘ��^���k�F�w��~�J�Cr}+�Jһ��� �dj�4<8��r��8<�X�'�P�1�h�ר;��gS�&�H"Ᏹ;]�H�?<h�
/7+M��҅a���d3Щj�oS�'4���oͺ׵N������?�K�<�r��`�`�����/@>�����z`I�kO)Iߓ%K�WW����SL���'�\���zZ�jMA�)��*�o[I48�""�®���S�;�q�r�n�s|^������!�
Lη����!�R��'�")+��Q�-VɠNP�����]�^��3�)���x1T����${,�ٞ� aa�Ֆcs�ǿEy��*�`pd*0�w��#i�<Zy�k��MV��^�(�z���T^���&���+N��J[�n�Q��G�C8*F,�z_�U,��iF��3/�R�n���A��Pa;П��L:�!7'������H0."f�ζ�(䱦�B��;��������h%�||o�Â��~2����(Ύ���1T��t�jW���d��H���1l'��@�@w<�u��L�
�d�y�!Y<}>��B�}0'Z�Oؕ�!�����ɨ�����mt�t��H�rS��E[��~��	��'�Gű-����G�k�]We��R;��ihRO@&�?��O�݌W���vsB������V���WFU�����֧�_���T-�,�KP&"�Ȃ�X����Ȥ��t�fpe"�C0�e� y=��n�S�J_��B�I=��(,s�12�5��}�팓A�F���47	��ңsҳ�eM�v��d�Yi�@k�	���R����r�C��|���7�L%�]s�=��O��e~�҅H�*훩0�w� �cQ�-��G���ʨL@"X�N-��v��j��U4�=��A�0��ME��	ď;��#׊�P��a=u��ҍ� �o��8��<�(�̓�l�e�fr��]�9�<�;6Q���s��ο���'��vLnQ�"`��;�W6�CjV�d�n���켢�gA�ߵ��ͅ��u�0�G��ic����t�-CQ�OP��kY�? 6���}5�wH�ByjY�Nn<�{-粚�s��x�2͂���D'm���j�Nt����4Y�o�	]�V��͹L�\qD y����H�'nt"N)�}V��pj��8�1Lue[�[�>��ɷ�n�	���&���[��1��+��//�o����[�%Á/ox�1WG����|�;P�c<gOn����ՂM&H����ap4�B�<
��[(�V���7�BVi�L ��^ ��sZ=���@<UL��R�$%��Gc>U��;t�x��M)Z�<�Ԑ9x�"#}��*���^�2�K��k�j85�!r���8�R�p˹�&K�!��J'�)�V#�]Yʍ1V�]�{B_�)ЏS$ս��ubo�娠��D=��i�v^\TӅR�;0_d�<����V��i$%�t�7���9G��ә����>�4���������ϋf�ÿ�:���:/7VkXRA�ݥ8/j��bk'l�����S�r����~�Cʯ��5a���̓]�Vj�*���;�J��&��F s���r+�=��cY'�h�t�i�ʓ��.���c퐿����0Z�d��4ӽ�l�+e�D��=�G���M��?�ŀϼj	>�a�ECl�l���i���m�y��ٺ�m���s�Pe��9�%��������g�oƵ�ǱZ0/�)� ��g��S���ŵ��	}?�r)�(���6=�����+�߇�Mm��TҥS偈�
��"��tNCO�1�7�e�e;����9Z����������=H�t� s�k��g�%�D��a��! �9�qp�_	�;��o^gn��aq3��?�+k0���#��YPN��O$�P����3�)$�:xk_��i��^��E�Dq 쳺 �`^�n��0�߻�?�DY������\)��ģĽ�K;ˉ���y�u�܊yQA�O�Dh
A"�~"�D��� Ix��2���0I;��(�O�ȳY�x2vǧ���A U`ɳ;޾�l���"j.���X�Pp�RW��.^3�hl}��_�|��~�w �X�=��Y��G����l��6�{^�<��\��VJL�l��#��G�#���Vvj��U�3_�].Ћ8��l*
A{�J-b��A��P��[�0~����2����+��2�(�c�/j!Qŧ���0k*�����!xLN��D�K�)?� �&�+L��� ��"t� =�^��3���:Y�U���@����1<!d���el��0�G2�M��z|����H�a�o[ਏ��G���1�,�莩�81��R`d;Q���"?�Y`�{�Ksz��t��:gʦDK�>��,������ ��QP�D׈p?���_Z��'�I���������<
4���z��-g{D@�p�����<ڿ�S՟�}��4��mÊ���g:-����#*�Dȼ�,�I�"��ר���p�8zE��n�C���.��)�t��[ٛ��=\@j
�&�8�*��C���qQ��ґ�X����o9�"�PB�:L&�� �w�3(�1�ǹ�(���'aJƿL�5�G�z:y�.q�������|��_2�ܢ͙���ҹ�&�r8������C�C�yr�Y�>*���i����9x�d^��<�;�tna��Ro�,�2���[�o��[R��M����sJ�2����>���J(�+���8���/NIF)n��,�����c�y�5��<�Kl��#B�:	4�%�xc�U���� ���O��O*oAJ%�6w/��\�`��l4V��I����{͸�!8豹�F����ʃ'y̜�?���EM��ց����j�@���pz=g[B�f��א2.)��P~��w�ӢyNy��o��T�o��n*lŊp�e8]y��~`���m|s��0��@Z(�sl_�֢� </�6��*�߽K(�Cg&c �'�5f�p-�O�]�j� ��}���f��Y��.;�Ͷ���U2����r�fF���l�Y�ֿ�k��=ѡx��؈�=:���T�b��43��*� �Hq�� 7yo�*��4�tvE'�U�͒}q�����7�F�ߦ������/ň}؆$y��0f�P���d$.'�3���Y�س2{0�ȹ:�誋V�g�W(���&��g�N��& ��;��ّ
G��̃�����pj@��<���{�q�LoQS�*q��E��y�#A2��=0�|{���p�M`��j�AB�	�D�V��>���ݔ��0G[�*l� `��0ڿVP�boIe8�!��&�KĚO3UDJ�rx׍�Bs\ӧ�(�Ωk�K�D��x�={�#��/N4���ܭV� ��t�O U�x&��T��/iӊˇ�)%�+�j���u!QL��d�b�i@/���8��F2F���L0�^�P;G�cm\f�ઠ�s�0K��s�<s���]{V�1H��	��9���!��^��7���� �"��/��} �MA���;LP����*m��p�/��ftӭ
��~�	�@Y���F9���H&�=&?�+�?���oBb�
�kI6ջ�"��;�i��|+�m{��UwwZ��J�L�-�Svx�&�� /%M���:��M~6t���>�3'��CS��9/��+U�$3�_��#��yN��&Zk=��u����V|Jç��kE�'�&�.M�"o����ܦ�
���x�����yU��8�,��%��$:�����Әw�T���WBㅹ��@^�m|�*V.�sG��� ��_�Twv�BȈͧ�
K-S�S��
w�{�]�k��Z���ǫ$Q4��G��c�t���-'��Bg�e�c%G�Y�p�\��s���n`��\#��k�"�l�~�ҺN�k	�����n�
�J>`��&B~�]C.�/����JXY+����zW��'�ӣ��}�v�>��TL5(;m=�[�F��
'=�&�r�I:]d]��l7��hu��,��%���춆 oeʖǖ���k}�Sɧ�B�c��X54 �:j.���[��U�א&����Z��7Jy�0���Ʉ���1K�*�`wJ^��v�Mމ��!d�nd�����7���n#^6�`��`�Y%�$\Z�}  Τ��K����U���1n���TAuA�i59)�q��/����������4<�3`����ڦI��v��E/9P��@|������:�̀$Da ��G�:v>�N G�(�s��z拰�YT��C��.o5��|�sC3GX1��5��M�D���S,J��aD:��Qd�����-���VCd$!A����>F���a\Z�I7	t��Ek9e57b1^������}O�����}F^�Xm�A��/W<�󒞔�S����Ǎ"U��84|�!�.�=�ˆ�����3Q�v'$'ʅ�|�Z�Iw78R��˅k�5k)��0�D$�
�Ն���ꨤa��G�!��[SP��'�(���g�ʏ���@�wVֵ/�g֎AN��T��WPt]'~���g6�G�,/6���_j�X���iZ觫����zal{�/���C��mƞ��
n"�j�\���\7	s�Ɠ{�$�p�kkK�V�n^W�Q	rbl�Gi�qe��xQSf�3J!%4�ѬR��*�����7p-�ǀxF�Z�"�e�)r��û�����ySO�Ki}��< J�١3s����K��1�A�b<��L\�,eB&%��������d���ugv���=��i����6�ۯ\��x��ɋ��F�ú�{��q��U�,~W�|���8Q�y[ow|1~�W!7N�8�#�|q�ܱ���O���ۋ���5�s�Q���x��p�
_?F}gK�2�P���A�0�c�<�>���������9���iR�T�2�`����?����W%����Wq?���C̿��{�8����:dq�������֔�x.(��g��	���ЈK�ƻ�a�+C��U�Ad�c��o�/σ�����@ԏ��a�^Z}� ����֎����V���=��&l�n��O��PV��hќ������<�/�#W}+�����|@��0��X+*90sΤ!�f
$>؟bґ����j�=X�1"��p'���/c�|���{����{� ߦ�N�&�h����x���%��}�T����b��V�F>�ݻ�W	��1���IRc�L$����0:&�m���R�n��B����Z�	�f�N��
��;�X�M= ��6
7A�x'�۸mˣ"��z�x���Hno�����ު=�<d�2��F&R���f��mCKP�L}�_/dSq��RR�lrnmD:��(3 ���LhFSz I���ɕ�����W'7G�죥'���-1���Aᤣ�O	�ŵ��@�v��m�L�zg�
L�{��?6�$����+g�+XUM����$.�A��7���d�
�.�٬����E��~89�E�;]{��Fiܳ2<[x�8]�%�������B��r�#�%���.�0x���x�J ��S��8�1�CheBy�Ut
e��0e�E�v+����y����=*�I�� 7���
�|���o�U��V���6$�Z
3�D?[DH�f�I�R�4����Q=�"t;,�'��U�9����.cr¬�@�rpd�j3ͦY��m�y��H��$��6�����'=豂l�|��N1�4�}_���bRQ Ju{Ճ:ra���.��5؋c�Ƃ�^�(�NS��Y'_]-�J'WB��ب/��Tk�K��1�*2@4�$ii�������狯���{� �(�\�H|cL9>u��֤�5���=�NX10H�UǠ¾6<ˇac��)c�8m��W���]�̮wb�uA%j)j�S�����$RzEɧ���4��&�;_�2^�d��f�����t�B����s�R�����6���7�����<�& Ug��f+-t�����"+���{����H��b��f�Ϡ��蘒ݶ>cF�d\�<N�L R�)�ЗA������8��O�ݟ�W����Ϣ��<(�q%-���~��8|���9l��TI��m7��R,��ve0O�1�;�V׌:"�IJ�y�U �{Ē6�m��ה&ң��9���؂�u9-lS�A����Ow�O�ܭ�S|=��]8����b&mM2��`����OƆ��WM����\���g$,`��͡�3or¿���&`I�T������@���4����ύ���m�Y��7�l��Ǿ���/[�X�1f*%���e*��D^�6�-j,��� ��p'��gtv�V�Ce.# ��q��u�T$�*�K���^ma�u
Ŭ�^m��_�ch�&K[甒/%L��1�,3/��ռHi�����/���~�7��u97 {,�����05$HT���	#uky�� ~�s&�K�(��`i���<ݝD�h�Dk�_M��H;+#NLNor�}�W���/���X.�O<�b������gF�tkʯ�q�،`����Q�����8��|w�űl
�=65f��`A9%nc��G3���`�7M�����0�N���D�ď�_!��Z-�����ʽ�,�����?-���b��Q�p�9������v����*b4ߛ�l@���!哞	���h��'X���Q���m��Η�Ʒ�6�eYҢ���6ʻ�3�K�U��[��H �����T0�%�Q�]�WP��Q�+�3�v�3kٿ|+�)^J�u��=d2��.�-?~�~r׀��6^W��Jg��9ha�h�즊�K�}�{Hs4�2�g�k���x�f�Mϧ�84F��rR��t9���%E�
Z�*�N\��o͌;��	N���S�Bn��|��di;G�"'k�"[��EG���x@H�'Uxr<��fQ+�l��GJ+"cƪ)����
9�tJx����l�9�M�%S=�&N�C�LD�iE��F�Y���+RN-Г�ة�$�P�6V�U��WZ~:�X�fðx��ia\p9cd�DZ�ӥ�ˠ2YBa����X*�#��J��w�����+0/]�5����l��n�Tŀ���HH��R�e��2Lc��_cQƫ&��o>b|	I��o��o��>u0��Au�Yn{��Ф��C����Lm��-yz�}D}Zڦq��:������<��?zG6�-�[%c�	��?7�<��^K�|ˤ�}.A�[ȫ�2�$2xW�]��ǵ�d�/ v/��p��t��9㖽Ɨ�P}y�^~7�B��,]���"̑1\'����Rڥs�pk�5�j�IR�/L�oХtM��pq�تà k�pcG1���1�evAv�1
���F(��K���!K�{�|�����K؞Ӡ��X�wZ0M,n����1�@SfIl];�����m<�HM-2w���ؠ]����N�ETOcb{^*�Y���� 6{�f\�u����0���i��y�p��c�)�����Gaʡ��������vL7a^qЃ��l��ƕc��z�o�H�h�Y��� _A���
�#���'�cU�������/�=��#·�f�%f!�?�>ﺭ�wx���>�3�v����uW�妩�Q�����(��\��z�DU�:em�wBSf=���Z8;{ȰK-�u�M�k�4��o�+��6�3�oT �|	�̊��<<M�?�����4�Rt�/�tG�7V򈉅�ң��DɀlG�`y����度��	���b�T)bf���z�f�ɑp_���w|f�򡺗� yQ<Pvq����,J+���g��i@Ӟ}I3��=�''�\��)=�WFÑ`�Ɇv~/o.Fp�YF�:��t:в���	�ހ�D��M1�g�֛��9����e��ztDX����{lD�j�V�l��Dh}�=���5�Ch�8�O([��Rd#j��b2ْ��K�ݱ������,^O��j_�]��)��qv	PfN>}��R�h�?����n���ȍ�Č(�;�(14�J��rHe�O	8=8���_ �4޳����p�m�$�A�iW�Z�����\׿�EG��$e�� �@�x�0s9Q(��q�Ɣ����ܯ"s'��9C�eh����U*2&�@q9�Bh�>�e�����k�g���X�}PۓL�tۂ�0��Z���c-	'p���F٨�n�eN�"���\�zݪ��7F�P�3�$�)���'�H�_�:J���1�'x��r�<���*t�(�y�@G~�氪��Jҩ{ke3er(k�US~ҐL��7��9�-|��K����y%շ�v%k*�0ʲ/�孚X���|���tڢ,��xrl��g�����q�g����\��^�#��Rơ3bn��(���8
7*+-�ZH�M?������;k�UR�Ki�28Z��t�����[��m������U��_L���(�7�^����8��ڪ	ҹ�[ֶ`��!�;�O���]x�-t�+z�ZQv�����1���@�����/���s�龑_�b�	#t�鞒y?�ؿ�܎p|�n�NO!�ה�IUH����Ƚ�Y���I[+i�'��q���_C�L3���iB�������tf���L�����R`���k���E��1�\&K;��e�c�;���"�+9a���2<[�J7�&��ʘ�ǹU� %[<yce]f�M �H"'���Q7�XxA��h�w�������P��HcĎEO
�FX;�{δ�����Dr(���'��&#����_��Jё����*m�~���Z�$?H�1��P��d��	|H��S�$;�,���ȱ�O��?$�`)c������tE?��qeМ{8 RJ��e��<��D[��{&^U�M����攘�;,�|��Xy'���;UP�j�
�ۀ�������b5tvH<���ߴn�h�p � ���)4⻷ݪg8���?���$�[_Z������wD;&ɭB,b:��rkݦ5�Q�	�E���hҶ��N�	��|��2�� �H�;?7����k݊�uW3��
� Nk����1�*����ʱ&�o_�����Tɴ+X�KFug{���ju�P9*��1<��x�	�Y?]|"��1������H_à���8#�>BU�Fn̾�w���5m���,F��~�����.g�P|8tV�3�B�<Z�(��Q�#�.��&�Btd�cW���*������p��#��U��Q-_�,��B�C&\cp�����_Ⱥ~hY���{�R����-�U�e�"�
ڱ�^<{HM���Yݵ�V�7�H�ў��o>�����Dh,(R!7#���b@���:����c�)���U�(�����+�+�5IA�,x�μ���.k{r�B8�]�d����v*�7�A4�&\�9���7Fg��/�����i �xN��nv6%�N�^<���B�*��RQW��V��4�c�2��>���qn���������h�K@t�1�ȴ� �*{�?��
%l���;�-y�-�Bٺ>�I�!}�-=_<S�ه4�؈Ї�}��`�㡊Pe	-̣vln޻/R� ���ߪ45r�
����N�*�\Mc�?R�$� ���A�ҫ�c��O�G��Q�q
 XCwʿ�:�x�e_�D4���.Q5l�T��Fn�5>�6�W.�Ka�"�͉��*���Pi�{�sP_˚�6��]�U��y��{��K���e�֫�s4U�*�=u�X*�'�ю/C�K&ţ_ d{�r�梮�:2kô(&��3�
��q�Е3	��ӴYj�S���@��J�P�����:u��Kd'A8�rYaR�W�p �~�3�`Y�j���'g-f���|T�H�;� �"Ӳ�y�V���Y��z_v�g��?q���+\^͈na$�&���ĉ��r@�J��2�[��(^ȍ���4��  ��.�Y%@R�+v ���B^bAZ.B�*��4�&W�2An��mhO�i�d#3j�*�S}�쑤�~.8F���`�(x8������Ӌ�^�җ��yMκ���fi|5�>�3]Җ�Xv����d�xot����<�Eo��,�i�k�$��P.ٛ|[r��"�.K8���o3M�Z����8:Ў�����y{��b�Qc���L	����;��V~Бn!D���n�U�1\|s���a�A����|��1��k����,C�'�Y��sa�����;�οA��18�8/�o�:��Ӌ!`h�p�tMQ@9G�>��{�Sb��Q�x�{�n�n���5�8&���@C�g�6�e��7!�ȇ}Q+������5�q�k�L�>e ,���<���b]��mfUN�dݯ�%�����Z�t�*}��H�>�o�ji�]f�$�{vi�,�|���Ï<����SW8}*TRd}��<��rM�/�Њ�`�k��j�f�(���e0wΣ��.BAx�q��)��	�He�*[_�t�����ES��8䉵�,/T��$'�t� ��T����ڼ�D���T�\bb2��t�?�P�<�^�䬔�ag�i��8�9q3z\b��h:[+�Pw����e[�+&���HLw��f}�W�M�h�M�ʒ��|�#4F�W\{&Xd�T�e��U��h���[=q� ���unc6�MH҆�nY͚��F!��I�?K�DHF���3yg�Vסȝ�}�DZ[׮��%z,)�Ϯ7z�E���W��L��K��� 	.�����n�k��p�e�虻���1+��p��|{����G�HRH	)ֳ̯�����$~��K��}[�\~�NDJ)�)����j�}�}�֟k����C[��d"-��N�g�1򚈴�}(�>����
!?Y��.D�*��{��M�Q
zu��#�o�%��j�s�lw��m_C0��;���b��������hE��/14�x�3˷#S6h5vȌȾZ�ᬥLv�[$��z�;��Q�2�����Uh$�h��_��J����9��"���7��I=��J�5������n�b{�'~���b��բ �t�c#��St1�ޠc���ʦ���U5I���:>&��K?Ĕe��O���m���Y�+��~���b�v�H.����O��ET2�Ȏl�l#N"N&�I�؝GS���_��k'��~�����#���7f�3fe����r*� �5�OֲP�O���ע���h=��}֪≥j3Q����F���z�z������,�u<{<��^əM&.�1�7;�.�BA��C�'a��
�sx�(���ZQΞ#7B�卭H �����H��VkǧÒaZ�Z�q��
E1(���id����ă���L������Rd�4`�-2b��_����0��ٳ:ܴP�zm�`ͭmW�~��Q�eȲ�H�T ����-<���LT��W'	��c;��~�c��[hD��.�KNo��v [�d(��7cG��λ��~�L�aB�('`H����&D�v��}���rz����t�Ӟ��ì썣ꔐe�7T+��)o�ݙ@K�:ܰR�H�Ƃ���P�}n5�ma=KE Ө�����4��pB.��A��DwzB��鯕���;��<���� ��5Gsz������	]�슽_�F�+.�h
9p94�4���jJK;P����.���v��;�=��4y2�b� :��KLi25o�� d|k�6 	��ԙ`���? �n6��� �e�yk����"�Ucc���F+�Mf�^A�B�y1VU���OR�7�_c?+�z[�ou�]�7�W���z]c�Pc�� -�i�� VU���&���ؠ��b�K����w�y]Mnњ�oQ���<�+}���3�N&�����[�gH���g9��"�$xw-�k����_�2Z��[��O�T!0B��0��mgoQPǗ����Jck!K�^
�,�=�E��/�Y�"tW���}��~TV�2[:z�����@��Pe�A����qJ/uH_��.�s�0��������xu�9����?�}���`=�5����m"�����];�(��p��
��پPu�s���cX�Wb��Ba�p�;+��=$s(�:��d�����C�n\'�1��K���>��n�m�A�T�S8��GW&5nU�-��̄KT���|��מ���
NE�]G8U6�^����:�/�|��[�6f��:^�V��	����-����2K�c���ac���r���=|B���3���1�,]��JZY���� 8O����?vY���wIT��SF-k���!�QA)'�@v-��x�J}LsC(#�m}�G�̞�R��6|X��"	�ݲ��W��u�������a�)}!��2K��ڜ�%f�6|�wr.%~��þ�~�φ@/��+����D����#r�	Bx�4y�Y��wIv�2w0
/������)��OI�r��m��ޏB���#���)��K����A"��/C���N}���'{��v
�6�������d�'" ��3���`�[.���v��T �	�֥����bVO��"��c+/D�8�S���� %]��n�-�ʠ�-��b�-�d�ؤ�.+m�<\p*Z[<��juT�L�睒\�[�nQ����1 j5T��� 	"l��qOʛ����-�E�6b�E:�ķ�ܐ3X��碽0��x�hf`�4��B��Gګ^�Vwkq��d��07B �j;t-j�='Qĺ��l�4���f���_�℔�U��v�!9�'܃���QR-�fZ��ɳ�^w>�V��Qz����{�ڑ�$كw��*�Z���Uz�ܭ���V/��酛�W|ZA���ז~�B�#~�߉G��� �����ïҖ3��o�n�9���v �Ԧ�֮4Ȇ�x="����-�d�}ri������6_�i�FFπh�[2��R-��7�h����B�8`'�V���_)zq���B�c�VR���*\��~1¹�E3�	80I8�H�����9E���u���Z�W���Q��WZJ~�ݳD.`�`�(��> �'� �.��|i([�2���Ӏ�Db��(���Qy�h}F�@sXP$"���ŏ-�O��鶌1��k���;��hË�ǀ����`�ߣ�1O��LӍ�"�G0e|B�m��ڬ�>�2d����*bc�~���FiۋR�@(LX�#s�k���j9u�M^�3��j^�*T:��"�$D8E3ܬB~[蘬)9�}#dM��㡺#���_���(E̢k����7��/�;�8�ZQ��M�lp�bxħ��!d��g�Xߠ8c!5/�p���ޝ�~ʋ�����y�(7W�U6����}�^;�"Po@uܜ�n��44Z/�CI��h���*:��A�]�C��F���c�,�x�ʦUHB&y����SU�
��c��2�ɬ<��M�O����y˳r:�5'W���pK����"�B�Ҵ��uP���PB]�Z�G����S���Yc5xK�`��Q�EX�L^�*�nGo`�M�IKo��,�����2#
#?�H4�����K!*���
��V 8_�Ձ��B��f���B�
�O%�9/�ة�#�܍�r=��2��VKJ�r	1+����KH�����w�˗�����J�g� r)��A��.��$G�wz�$~,�.D kW������٧��P��P�_�FCT��S�n_i���ڦ4ǎp�n�⹚U���`|���v|˞�q�^c���Tc|~Nm}$�wQ�J��TX�:�>�er��Y�_�H]H���)0p4]�<��o'#��ş�V(��ipvH4E��Zi���6��-�;�,���& ��/Y�#�M(�v�s�����ɛ��0uQ���A�����8�X*�wjc0�y*A�TT����,_NE���._��׸��]'U�yシ�\���L��r��ы�ia���xPg���k��B^�E�g�tԩ��������kwx�Q'�\E�i�ك��v0��{F����Ӕ)��Ւ]1�#�v@~W��n_�$����s�^�4DD�Df1!��E牐��@���f�-�dR2��	wq&w0��[��CTa�������z��;,<^���Z,5��������uU�\S4g����M��>���Jl~��
�3Q�\~��u�	�ɔ�e��!L����G�ȭ��d1W�~���Oԗן���������B�{,Ⱥ�ԧ�"��T���ňL/re�����Vd�x;�դq�O]���Ze�(gO��@sU}�q_�A�ȣ����o@�W�"#5Ր?.�4�>���X ��5���Q�F`N�����l?�l���ثm�I��	+�/���!�C�vH��A�`|\((�F���LƁ����v_��ا��Lx�Z�?� �ɦal�r���̌O�V�[�E�����w�izNQx�rpsC��܉�wQG��Ϡ�4�ȁ0�����2!���5�4�ȉQ]	_�!��a�ތ��?vY�kҼ{�8>�\{s��62���A⏘1��� ]K�M�`@�v�����0�����^n������T	����q��'� &��a˔7��B�h�dxy�m�d2
�ӏ�e�D�ڜv������H��<��Y/u�J�+�K�o��d���랴��:�=�B��N�t���"���8�bm|�k�u��r�s�2k��XDw�eL;�3=���:ڗ&��W߽��W��2�r��S�v��v��:vn����Y������a��=�H ��]���I}�!����ЕnZI:�{ׁ.x����6�R�OԜl'e:�I�:���}�Z�*�8�b�Q��@ŏ�]�T�tZ�af���_
U �O�M~_if�4G-J��$,~��Kҡ%��1�8�ϼA��$�y!�Q��vW��}G��׳q�צ~ݬOR���`@Xm3~�M������N�I�u5�1�����6��ڡ�rd���hFh����4߼�U#���N��4�����)�wljj��_)4c��i�� ��iF�m�QҊ���/��Q �Ҽ��`�����sБ8�jY�*� f]t�Oc�������i����
#FJH�W�=����S�P�r!(:�5��h�-ӛ��>Ze�<��K����*�s[*�-!��w�=E0�D�����Y�`��'"�}��y�^�����fO��HT�?&=�#�uc��9�ɘ�Att�����#��~|)v�]�rm����|굓:��`�?�gH��K��62���CT�L�b&)�_���;et9o"�rU�ޅE`��5��س�"��X,ef�7?櫙�_�K����kV,��5����V�5�M??j��0���<�^U<���
��C>� ��-Y�U�W�������S;?\��0ǣ���Y�X1�	,]����O�y��[չԔH���s��>�JE��hI�����+��V�����:�sgWa���$~��K�%�����c��;�j~E7m��n4���Z�~cJ�!���
��@ly���&�J}Z���F��J<��7�J���0��՟Պ���&��#�<m̀6�E�Z�������m�e�zZq�6�X�-��]�=�*EL�?�@�`z{`9�Z��eƞ���Aa��2W����z�'���:��DE�9��Y 1�·=����c�gr7���,�,�UNdϻL����U���!��o�j���#�~�IbP�NR�U�c�X|��; &q(��[0D�p�`	�5�/�{�>�ԙF=O���Ѱ��n�'H�)�$�|0����l<3�0�b8����`P�
*�Z�����h��̇�²�y�+$����|��nc;�o:�����
�3h��4`6b��2h�rHM���bsu^V�b�v^G��:�`�j:o�=v|��4��s��?��i�X�X�ֵ�	v�&�;V�Z�g����d��==��?�7���0�Wę����Y�f�6szGA�2�eO���;擝q����Z�,C�#��t�z�_t�4������)J�Hh�q������ޏE��#w�e!uD	��9~�I&.y���ˁ��!��:n����X�iI^��\S��]0��B>� !�a-u׿�4c�-��v�.��v�Y��όֺ/HS�Go]�ٟ%�)�����-[>8��R����o[��K��T$|��ɘ:7j~owpkp���x���7�b�������N�������
/Z��{��#@�X�Zv^�X��*�!���]�?<z�,��MT��R��{�AHt(t����;y��Qs1��.W�)�C��������fbRz>P�@ב��m�X�G$ dS�~�b�H抽$��H@�N�ƣ��L}�J6*1\�4*��᩻黵�k�E�1.��8�ܛ�Ԫ3���0f��(35WF�G4B��(�_�uЌl����-/ $�O�,��Ӹw����j�����d�+Sh`~�e�"��u_��a��#/�ུD�X�!m�_� 6���n�Sey��he�����%w{O�&��ŵր���r���2��� �	F�[b܀|�98���w�j�v�����y�������Nh�>Bi&�=�I"x�*��e�%#�/��1�H��K��yehL"#Â��{⎥ͣ��F	�z0��H2*��6�;���]�ז*�@��Y����Rx��&�C�}&��X����F�&[Ѣ�9�\I1{�����^'���~e@�<��p� ��Bz����r��UP1f	��POڹ��$�!���ZQ��L�0��4/��愛
���}¯~�#�)�����w���B�%�)��B�s�v-���B�(w��0j�x�!5�p/�l;66����%�j Ζ�Mf?g� }������*� ���Q����^S��-!��cu�4�Iïo
�1QH�
��Ϝ��Ğ(�h����b�5���Ŝ��h�8�L*���e9�h�L)zmq1�{z���Ljj4Zṫ��"ж�ef=�؂��Nk/��#`J�kɓ���5gB�������*��2�y��mS=��_��[����Yh ���}����>]�q�����}�Ϟe�f�lv�yTxU7�?��P~V71�f]�ٚ��f��T�����<UșuQy�֕Eˣ,��C,�6!^�H=�"����+?Pّ�cb��Yj��q�J���ʗ̆��c��^~�t��Ϣ�vuC���0Q�G�؟l�_�兼�������+��m���D�����[��,�� t��ю�J���q�+OH�.Y�ў�mk_��U��>����M|�M�{^j7z�{�}�9A4���̘v��kaz1�hg�A��|F�\����\�|TH&�!z�󿜈C����ne�?hN�f�Ih�����`�/��O�Z��TTt(���O�Eo|��7̸�}K0"0xJp����e��\.�]Mc�t�f�A�/�����E4-l骂o�#E�]���kTV&�]�(�1սc��w9�;�[Rx���:�ژA#�7Z� -��r<�ҝ���K�0���6$��|���� M��*��V���P5.w�e�Ն�z�|�����
����� L���P�Ie�������Ih��i��f��� ]3���P�o�4?_���� �#�eĆ��ڍ]��R1�E�a�|7?gG�t��3`#�@^�z4J��Xa�tp��>��g0Z���Hнy:&���,a&�b@��٬�?�p��p��~���;U�1u�^��ͽ���L$u��#�b]d����aTv>v�9�Bjl�f�k�O���FS���ϙl�/V�H���5[h��9њ	"B�"X;X�}D�f�0�B1��,�����,��z�Ӆ	����!��� �e�T^D^)S祖���Lۥ�Lp�H>옟����
��h���BQ)���w#�j���H�n��R\�٧bPl����	���Q8��6}|���7OIx&G泾�_H��"D��N�as�����SRA����ٽ|��1v�+���	���nXG�?���!�39L�T/*����zh�����8TH����K�,IL�0�xZ�����$v7
�t���Q�r�¯{=�Q����r�m*s]~Y@�,o��eq��>�Z��o��&�8"�R�m��/�ڍ�Ck��s�_���9��.��Ƃ�"�Y���3 1L��3����ʹC�#��w��+H*\�%9$��h�S�H��W;���Π,��Kq$Ak��p�p�����!-懢���r���f�xK�L�m��娲/r�ѰĈ/*�翑`��#!n4�~�%�;GW�"9?��	P�L8q;�-C����>�z������@��$f�$6�=�pB��l*�X�����Z��Y��a��`7��W: ��Rz���Q5Z5H�k*��gZ������̟xE�L,X���͹;�A���/�s(_��_ɭ��i*�
�nP眱����0ޣa�:UR+����(�qS}lŮ	��=�Y��@�b�����c�|���ifЧ]���4���+/LxU������)dhA��k�Qת�3�w#;�~u5]S6ũ��=�o��΢X\%�$?�,8�ާ�slH�U����DFD=Q��z�C���1/Y5dX�]�ߪ��u�}$��B��"�R����$������Ы�S��h�I�MT�Y�^3��M�J���a��I��u땥�Xœ�i!�N{`g���p��z�a�{i}��R	�aG�C���Lrz��U da �x��-į�+�i-Xv)��.�{�rø�a^������FV�\�І܃T�0�]�@�.�?ѥ���tm޳��X8s��D�=+���#'k�8c��.:(�{�,�c+b����������k�n�V���kРt�M���r����)�y�����k�M���qu�O���
#plK��/�a<�G��B�W��T�OE���.OI~V��FUes� Y�W��U�h|�N�1"�$�`�'\���,kE5��U���X��7N���`�/�8]$������dUO��F��u���RH�����Y�*��������ͅQ+�gUVi�k|�p�p�J�Zڡ�6��{s=$��c�=P|�N���E�`�ZS;�B�be��glx���|�'&%��+�,2���ئP������ go?ˤ�Yd��##2꠵K����h)�S\�/��P�}�l]���T���fkv/�!��TH� "�^W�N�������(\8�i��qH�&���|��t�>����[gڄ��j���E��CC7�.���ﾖb��n\�6s����cZ��f0cE�y�J��g�"�m<̀�X���INXX2���"�\�u���M_�ա���,��x�O!�|L~��'���ڨ �?N&��?W��|��`��o�U��McZ!�";cS�&edR��x����V���~;��|�gڋ�+M�9���u&<�ge��>G�M/��t+�1�uĳ�܇4	��(�V�hO�ȓúU��I�.���7k�柬'�}f�٘6��|�m��"P�D��N��H �T32GTU�&�!��=nX	�O�Q�bP<�l��!�]i_dP�q$Mᧆ4D�2+�� mL�7��#��N�I����^M;�L����訢����p ���rb �h&�\���I��0n7�^�pQXAx�l��hi�X�w]��3�ηɴ}���e*��F�<�#�Ù�(�[��!��JY���j- *}
�1O �y3o��6�ω��K ��	;��1{��2Bk��j��$�_���I��߉�(ސ����.{`��ۻqrt��-Ů�Z��ܚ
�$m��#��YQ�n���������.xm��
���������H��o�f��LG�	w�/x���u�c�UdUB�@6�-�F�Er銿���.��>�F�y^�H5;eX�h���\�q�SЅCS�B�u���q������A�j��
��/�J�5i��P���u�푉�6.ۨ���{��k���/G��a���0���@�*�Q7�mF�
�x���g�sn{Q�2�c14P�?/`�;�m��nb�EB����3e�6�
\���Ǖ. ����t���j2"@�f�RQ���˝��^�g8�3q!�d3 "`![簇�d��,�!��:1R貅-�����e��8�Ȭ��t�T�H[�!'^;˗�?R8��?�Ov�EO��Fᗔ�	Ha��M���������̘��w�uTKXL��5�b�f�5��I-�5���L�罪���v,H�pE���<��\l�ܸ���o^���:�)4�`ǻ� ���c���8o���²!�:ө|bk��>�OMz�^�K��i�1��;oǐ�Ȟ?
,r?�TS�C��l�ލ�H�Z� 2;��r�"�?8Is5Jj34i!��O�q��p�| �l�	].8�R����Uw����i���J�_�/�8��6d�;��G���"0��}��
4�֓^_�P Gq6��(�D(/m�u�����i8I&��ڙ��-�s��u���ʑk�S޹>i���K��p:���0�Q^��<d���0�W:eH�Ćכ�ˬ����b`�,)q���Ȫ�5��J#ʓT����1��!Өvl�`�� �l�4 ��w�֙i �R���PeOM��f!8=�1v t�!��;XBW���t�յ�p�}�=szW[E���q�.�ؾ�\~C���4˘�]�ê�������|���X�W#��*�����U�i��'�es ������� ��,:p���8)9CuU�D^RC��������A��G�9�<�o�z��@�2 6<��HM�,�Ǝ�Xfb��G���x��
�v(���~{q*�7�����|������ZH�ۃn��A�q=Cݒ��s6��o���H�(����&�ڼ�6�_A��y�Y��Z�XMF�,#��0An�(����@�;���j�Q�#N�/ᒼ�i�R0�A.:�\t�et�`D5���ekuJ}��xj8F�п� !9$FGge�6��)p���G�#�w!�V���L4%���B#�
���y;�D� �LYY<g���w�f�ɔ/�C��N�F2Hd��y)����w��J�����WA�㹅<����;[쟌"�s�b�ZC'�ߘri]c��=\��O�8Wp�	��V�F��tKKk3{�I9}9ad�ps`�Ⱥ���Y|3�G�n��E�/��M�q�ŝϺ|t�� ���A.z`�r�x�_~G��*��oĲ)YL�b�7���_6���d�Y�~'�E�����s�6AЮ��]�����Q���ՊѲu�ɫ�j�(Y	����������Z˪��	���R�\�u�u��Xb�5�E^�=OH�����z��+��BI�_�~�����Ɇ���wS�F�z�1�0|a�|�,u[z��k�T��ۂ03C~�i�&C{��y�x0��Q��t�v$���\�pωQ��$��g�$4}�c�o�"X����*�a��� ֜]z�9�A`�#�.-J_��BE�Vۘ��+X��;�O��?]����c����mf��}C���j�NI��b��_��������".@6р1^�`�%txa\<�g$��p%C�T�� �
$TF�������+>2^D}�\���<� 
̽hX�bwj���"qR?�:�8�92q�aWQ�s�+ץ�ܞ�>�"*����S�,��c�$��u��QQ��p��ՙ����v��K����0B�cA���Kv��ww݀�o`�մ����8������٠�VSzXs�n��h�74I>�mF-��/b�&��\�(`��\)���ͭ�N�e�1h�0;�ݞǎ�x>�m���Y2�JV�����y������e4��ۇ�1�P����>d���J���K��+u��wS��:��[�}��uX2	�\=q>_z�F_G�6:w�������9�]V����3ӡ'�������<�!��,:�Ж�'���өg���=���Kǀ���Lg ���9���m{��(M��Ԧ��&M�2 �۳�!D�h����-���i����}`8�l}��8�+g>���p�F���>io�;ؼT�۵�*�����o>�LgDF'9���щ��H��}���yፕ��u	Ag(�#���5��a��O�c��Ex�L�i�c�>�� /�c1���˂B�Hވ:Z�d觗��f"Qg�|��� M�ރ8w�%�+���/^�6��Si6_ �C��l[�eQ�J��
��I���2:����b��hnOw��BC�者=���-���RP�d)��� V�H� �(z�t��A����g�%����)6�3���֢_Ei��'޽!9BM�J�����jί^ΏU��	(DBz/��(O�y�RJٷ�����#(�����=�.�*!,2S>�>'E8C�(�{R϶��g<]E���b�����3_����Zg�f�)/���ò��]1%%�(��ϛI=���,�ٹ��2NG���ռ��zr��[
y�Q5�r/{l��qⅮ�����u)��ձϟ��>F��+�P!u��w��tV)�Hgu�訦�]5����a$ ��U��u��
�����}��L.)D4^�E�wQ�{��@�&�E���R�Z����Ӷ�X�h�x<�ǂ��D�ꮲ��+�ET�(3�Ω�2
X��I��9It>�X1�fnOo�ky����K���h����&!Lx��D|vb@�D	�\��?��9�α�*�'���4�s~��C�o�ݱʽ,��wM�ɥ�����l������m�e��`jOA����l�$�4ǿt�r��Z�e�R�W�*_6�2�sߐ��=���:_�ÔU��N���bG@Ĵ΋.[\�l�oX9�HLލM���J������@����}�:'����puKL]ɽ����/�Z��$&;{�{vw�9U�m�K!ԈŵX�Z����2y�Iq"]4��_�^pg q8GI�آ�pe<>��pU�@��ُt�E���|mZ���F�@�о0����l��OLj��R�qg'��|�ފ�t��w��>~����AU�ZI�᠖� Nb�ЍB���I[$��0�!����n8V�VV����S�m+��4*j��n�}U9u�4j(C�}��<�;B�xl=Ǟ�X���� [��iFr3���ޙE���L�E��$�Ø��X.|��pf��D��+�cE\?��@Q�٪�	�1�1���h =���G��g������c�%��-$
�9N�֍�qvq*������6n�Ŧa���i`�9���=q�΃�C,�n�ۚ�x�)�铠��ە�h�*!��!]�sUBj� �ݵ�4f��gNǯ���p��i�[ҋ	s�b	sR`�S�c6�cS�����^�S:mS�4׳��̲�B�X3+��^U|ޟ��<Z۞�)���Z�5��-�~yy݄��fo��)J���#�!���D�o^JT���l���V;�f\S^��;���Ŧy�g�_�$J+��+Znvm9KvC@�=�wu��0𨦣V����H^g�����z�`���<s�Ǯ�,���<��U�������þ�[z��Ƣ����`;+��A�+0s|/|�)�;LŨ�m
�Ne���1���C��X>��џ%�085�	���:�8#�o� 4m�'w�}��f.��:A��^*4X:��>�Ɍ�y0�����4������n��h. z�������8����| /?`_v0w�w�L�����}������򠶜��>��<k�)jV�����Rõ2D��h�LQո|��o����{V4n�{k�����(�Y����}!�96~g���0�B�.����&�I�?�>@��Ck�(��-����6��X��� 	�td��B�����'at�Q�+!��lc��'���Bu�-�mF�C�*�l��G�X2�\_0h).O	�c�/�Ա'=� �h�{�M����J�v� 7h���zo}�:^�Ax)Uk�F;�G�o��ɮ�����Ǆ=�*�E���u,�8��{0��K_�͎��I�_t&o�x/&r��L��,�I��E{��I��MH����n�	;�7�������N=K�ib�	�X;*1�ߪQ� 5�P.>�!b�y��瘳q���!	��0�#ň	u�ӟ�x�l(� ��K��oV�+���ᱫ;�38��H!㕴ɻ�R�9n�����T�IJ4)۝�+ط�Ov����X���7�}�.���K��3Cb]K�0�����0�@������vɡXV���@Fb=�����=F�:D�1�*�r�4X��9,S[t�����E�����齱�"Rgq֟�;<~��Dpx|r�x��x�Q��;���F��9�͍3�$vڪ'����	xѷ�V�I�!{�D:� y�p���b*��{�b��F�B�@wYFi|:a#�# �'�d��ovm$�`����ⰕH�^l���K�U0_ۃm�૟��h�����b��-/o�V�nACN����#6_���6�Z��Od��qΰI�#@߮H��d���� T
��hf��	jS/��E��S=����n�{듣�dFO��ϟ[�����d�=��㧝Y	p��=�����aT-�L%��������A��|����cm��dДGv1��vĤ�����Ԣp�}����(;2/�;���G��OTE`ӈ`���x�S*�ľ�� 01�;l1 e��&�`N"ߚ����_]Խ?b���+�b�G�d�nOޢ¡���7�d�҈���e�7��8y��ɋJ�Z�g�B�]��󯛓7T �-��Lg��yN#�������5L�u�B;R�Ek�;���.�Z�9��I�[%��Z(7_�G�;\�C=Fx��t�xܢ- �G�{�;�c�_��4�u��O��n��\������B��d� �Ҟ!W^;j�yV�M��Ce��߀F�������g#@q����5����6����虘	x��%9t�d:A��������Y�m�0?h9p�)�2������lH����ި�$�qa��{�B����{w�C��;jk�]^h)[�3-u.m�Ou�X>�n��G�,�{�09v��4�5����Wq��a��Cċ7�9Q! )�1 ���Av��	ld��k������=/�ےF�n�fj�h�
K)��쏷Dv���pMUlN�6��	��.�Z�L���?ǈ���H��{�H96���>�S�Bl��w�
גGj��nz1��`��������������A EpM��ɘ�j�����%q����{��J>��|���`ݕ-H��5��О�I�[><����nmDUI�]upk��}\�Ef��ߝ7��q��g��ĲIv���#a�ہWd,������ߘӸp�oǜ�[ɯk[rEf�JjZ�`�rku3��َ¤�Gt��_���Y+*�u�Sϋ�@�MB;z�M�L���\����V(����ή�Q�S�^�Ѐ$Dԇ�^"�U4A@Ft�bK螫���/����Ye�����S��ljeZ~�>_��}�\M��(T��pۖ4i��/_XH)b���
y�cH&�.�خ�+&�'���;D�82�4��gf�h�/���j�lg´V�i��/�>��|n�RmOc =
�c:��7�<�UG��\T85Y�("C���>^�\�6�������ܒ5G�?oŇ�)���j{��ȯE*�����.��~�W<��u��j�	�2)��R>��@��H�QKl]Ԗ#���E ��W*�򲽵�Mw�!A��$of#Ai�T6�uڔ r]1�ze�F3e��s3������ �,Ȣx��ǡt/�y��$���٦�j��H���r�DNՏ�'>��
ꨐ�9vQO��Y��s�	G�*���xg�Z\tk39'SH�wZ�s�?y�%(��;�ѳO�ߓ��I�Ԑ��9���?]�< �P݁сQ�?O��A7��Ł8m���U��h�@�Q��`eg��c��mЫwř��u^�̖�����^��pacOF>L�J�M�ՙ���0���!oh�;�T0�u������Db�84cJ(�i<�{,e�3�g��u�
��^^���]Ϳ�U����B1z�t�-3�����X<5��%(��\��>�>���-	�;b��*�l�U.������Q ��5]�(,�ԕy˺�I�X��qE�7�-�c���,�of\�Kw��~�I�\y���Lo7����L���#ْł��RY�����o�C:�`~�av��P�h� uQ�w�z��x6�Ec2�͒ �� #��'�b�T�k�t��)~nRh�쐈Lq�fc� �5��#B,��<'W$�/,�IL+�c|,犢�\�\��qDfa�g��V_hg;����*I>V܏{�1�O8�k�9��)�D�h4�㰏{X�i
�s�Q����7���dQ��DD����*x�!5�����s#��>��@
jc���.����&m�;܊�����Q{���[Qx��h�.�b� �s��bdY8�B
�����/��eWva���j$�($G��(�m ����? T�7"��Y��38
�>���h��9��,�cx���%l�k�	��LY\ *.bIm�<�8�~�(��Dӕ>��܃ʁi���>��j6m: ��Qd)}�v�A!��x������R7��u�r��3����-�W�מj�,7���)fX���u�gKو��2:��R���p(H�������?���O�A�]�ֹ���-�c���m�nͅ`�q]|9`'�#�x��Uy�+��T�ZV��¿�+��r�/3�m�_���K���Bj���Fq�m/Ń&�I�+K3��5���q$=�@$����է�f�=(��gf����/q%�{ց�n��_KA"ٲA�ˍ�c���]�2��w�~У��MD�#��}M��X�h���$NW������d�mR��h�6)�#ˢq"��Dh�B��v� �q[a[͊9Sv�\JEh���K ��J}l��`߃
�V�K���L���8��� ��z͇�oN@$��,��n=�gK��l	�7�d��&�_�+�\�*�藘�L��>u����7�X������5�������J
@�f��l�}��{�G�5������}�47,2��%��`{�p�-�v�5�L�QȈ�ˑ
[�ގ�����z(�^"�T�k{���4��>��F�	�����Ya� ��IQ9�Z:Lǿ���N0�̦U�SaR�ƺc�R�P5�48�<�x��3��x���\s%A��e�OT��P�C`#S&h�|�`eF�3�UOAm����=)b��'��/ ��e�~n75��/�_X�.���}V�!b�t�@G-9�ϱ�rnb
�1����y��#�Nc݁A�_m$,LQۉ|��X[A'���� �,�\$��m�q��f2�����bQ�H'��S�e#k��E�z��P%��4�)���kO[����Olt��'��Փ#]�yՇ+x{9X#Rq����d��^Tq���n�ƛ�Kj�҈��r��Q���\/A`NȀ���?����$���,��V��L@���<�4�K``��*�_t]�éM�����r!4���`a�zp�����6�J�q�e|�,w��:�s��4ہP��Ay�7��`��JI�M�4-2s6���`�
 �^���"Y�X��|�LJ�~f]���q#D��_��$�]l1�^��[�}�#h������R8���?�<���MJ�n����C�����&cw�x�l����oi���I`�2��x��Hơ@���&Xi�P�h,)A$�F�Y������������|����HS�߭_h�É�]�K���m��ɡ!�?
8��(���lc����m�,0��R<9����/'�'���z�Z�H��y��)���-�ř�|��1�K\�mD�gyh�����{���A��[�O��A���=L��: ���U��w;�0G�0\��i#�/�H0j�T����pqaTZ�Tv���w�F?��!<(kx�ԙr�J��q �,��	����e���e��!!���ɪ6q�u$�s3G�)�������Yٕ6���7����]<�F-$���6"���x��u�R�v%�.�z�T4�sҩ%|y�Z��9����9c;}��;�sC���ӗ�ȋXe��B�ȩ6e̕bŬ�ؠ5~
.���θN��~�1UY6�6���OΘCb�Ϫ%|�nڬ(��7~�t�ފٻ�tٶ�ߔĴ(���@�H�E����۸��P� �t��*�~3�&�/�h��/��E��_���w�.���0�dt��%ܘ�Uy�(�B*͑$@=INvB���	
t�w�図&6�TV[�i���Qb�4�X6�I�������y�9o�	��B���ʹXaPZ�d�+�8E�!Z�m+�d���8�J�Y2�Ȩ���mN݂G�\�m�
o5�h������C#��������ƃzWH�x��h)t���̤#o��0����;�0����������7@r�Vg!�TO��6׶����C�DFcLBU�y�T��|C8ۻ���Xc��\�0���6$q�i�6����9�#k��J���H*�[��Eô'a��`��h��)}��o���֎zr�'��l��Si�>C�����J��s0W�n0mhE_U�֖��P/oޜ��Gn�5��o�i�!mo�^\�2؃0V�ع&�M�g�/�T1��HLUc�䧰�q駅Ug��3��	M��n��q:�x*-^[hٽM���6�K���j�:?��ݙ{w�D�w�P�9g�s�a#R�$ğ7f4:��e����'2|Y�ޠ��Yn1��S�٭/�bB���mRw��"�C�b'���ڵ�tVL�GDU���L$h�ېph�.����c,���}�6����U�_h��^}�J����>LUp'5iY�J�F��6�Ҝ@a��ٗ��[Hm"T�i�i��L��M'}� �1m�8���a�_�Q0�[�Ԯ�3T���{.�_	�G�D��x.�s��J�qqa����Z��Y�i��fʽ������O�BFu=<돨�����89�x�90S�^<k$�����/{��Ǉ�X��UJ|�7����G�4]����@a�8������-l�1�j�~j'@����9�<
S�R݇�1>kd�v�Ao.(���q%c�L~2�PY��5��6�X]Cy@*HH�J�� �3a�ov��!���<A��`4t��?�DU=�&eg�!"*�G��e!����v��ܤ����m% �X�q0�=����J���Z���x�W�Z��*�d�W�j� b�|Ea��q�}>�\'��p��OAmT��l��9�k��:�����@K�]Ɨ̋�Z�*�^qܑwבf�N1���?7-�Kxz1��^6�O�oq`�0�X�E�x�5�,	.��^��t.lx3V�+�_����-wl���+��ε���F��a0�����˟]�S��I�VNcc� h�����N�U�wo����)���HWurR9'nI�#�ǀǯ�����*����N�;%>8���ǽ꿡N��R�y��˳�!��wj�
�=zL9��X~Pgex��U#��;?aF捖��Pu��4ǐJ-�e��BLI�1��>qW�Fy�N�6�EeL���΋�}�@~�2����^�6k��n�f
����n��<	���Y�HYb�=�٧�ܺ ̥�,��<%���	��G%����t3,�Ӥz¬���`2&�ry��Ny�N�7�������ձ��%��&~��b�f6ŗ����p�R�W�~��{<b�h�*y��x��3�B���t��-�[�:���y�)!�[�&?��YD��Ox^G2��Z��ez���`���o�.ŭ�!i}J�TҙZ�v�? �~�gGD�
D}_pZ�M��L�a���`1$7Iz�}�	)]
!��;*nU�RU��N^�0�\R7�C��5|����� �b��� j y���`~F`b�t���y��H��~�O���x�>1�G�� (������	dT�y���:U?�IfưLC�So���;=�ힶpA�e�k�(��ʆ�=E��F���r�|�-U0�����D���( ��(l:�9��,��UT���Kכ۲�����AKǦqdb���,�[n�cܘEZ���܀��{�o��ku�G4�$��E�F)z��=��7�G7�'�0�h���}w�����d�>��-X0?���� � l�bNÄ�~�x������'?�E��퐲$£�3� )�:'�4�/1+L�@��ul�^d�T���4ڊ ��,d�MDޛJ��(�Q��j��WT��� v�$<{�E���sn��^O򶧢 L:A_��"�Қ_JU��)P��ZV7[ɕ��'v���w��]��O��	M��O������Kʞɬ&�GX1�:�=��YLf�1�.�)Y���u�;V��<�jQ	�?d�'gLIl�� O�-̄F�{�,K|;�p�@��{��0㏠�mvo��T	�:k��r�gH��d}\�Om� +�!w@��˯,��gwR��V����ȑ#$����mA!��
�� mA.p�#�R0T(t��Ri�Y�ؗV݆؍�F1���?�S�~����r���5>�������kw͝[�&�궶8$��]�?7s�����g�He��{q�In����I&��@�ps�>�c}2�%x;C�������4F��?MѰ���n��Ɉ�M1���<|�ԃ�YC`k���z⟗��zTZ0;���`C{�mdJ�d�{�Ԛ�u�5*M����P~�El,�(#������7*
�����O����tfY&U
���@�y�(�J�Ϻ盧�[�x�D�Zaw��h�S��0���6#�9;OL羟��$\��2POD��/�q�La�	�_�	c��)�K�F�9 �z#�j����s�}M��~�:�iZ�����^L�6�1{��cA�f�B	t�_�m	{o,Z��PR�H��KWf�s�>P�"�&3�ՠ*��{��a�2(_��kN�[��/.�0c����`깊�+`eg�G��H�n��kf[�z�^�#���j�A|��C��V�Fz>SH�+25.ϋl�W�&Du��e��y�Y.�\B������TO��D�+��8W��$�b̦N�p��'8��b�!Ï��������pT����
3�g��gy#�H�^7V�?�.T�a/t{^� �ִ�fd�~��M�D̟���쮈Y@�￘J�:�f<H�F\���r��t�N��D�e�~S������t�Λ��\)G[�{���Dq�N���z�f�n}q`!�ӯ����_��\(zS1 �F���n.v�w\;vf�M$A@V}ދ1�*���^����LS�gZ�<�r�_�=��-)�Cvq�+���u9
}�e��7Ak9�,�`�b{6=�}��f�rHJ�����ٰ�g@����Kj�%L��P��gf�x�8��+r��zԪ���c�� �v�����"5������w$k����f6��s����+��2�ñ�F?h�b0X �"m�lJ�&��g�/X�_�p�p�P�ݱST@4J_����#���D͏��`X�,d��	"�H���q����ދ✼U����S�BC�Ҟq�&8�tB?�U^_O��rB}� Z�2�?���|�WN�o���W`����8�����!S����rŞ�!/�ӧF�|%�4|����1��~]F��B<�"��t��ug�>_����5|$ ���@���6�Z�p�S�\}����V�gR[Pij�U*�.47q�
It ��_����R�v	K�s'3��I��eF���q�Lh,W�ZD[� {9I�m�x���x���^iה]ud��``J�v%��~�N v$z���9��F�2q�AN������!��Y�O��Ӯ�d��3
���>��9b��pꖖ����������A��͝-QӘo�$�z���y	��E�AS��f���}P��..(���W�YBC��et˫�V�l���PS#T�)��\[��E �G�w�)��~�kTox=���5�NIP�dRU~�������iG��Y�ms[��]�����������,�� ��*_z;.� ��Lm	(�D��io����~��<s�X����
&W`�yۡݩNg���Z�2�NB�'�Eq�d�`&L�Q���
$W^�Yn���B\��ߵo|�3Q�URH^�(����l~��3:�+i������	>
��m9c���_M)QIh%��(?�<��ݲ!20�c���z���:�P{<�(�������(� w�w:*=��@�+�ad�@p[�kmz�����=4f��`��ٗT̟`Y�P����YB�gi�Ѭ��Ro���?���It�G+��4�}(���]~��WH���Pc%/��Ĵ�|�/�@��[*88��ɑDq8�:o����~'Y��Ҟw���C�"|ĝ*�SW�'l 2�@�:- �Nd��,;Rc�B���d�Ow�J{���؇�j-ę��L$�Ǝs�pW���s�=�֡�?Y4&~���뭢7��O��21�[�4�yX��%�U� �z] �˴g��T�0Y��������?I��-©4ǉ��%[ە����CxP�om~�@��n�6\M��D��zG7���]u�mv�
o��	�1�d@����c�V�b7F1t�I��A-�Sݣb�[�Ѯ�޸���!��;UC����#���Q��{�6)��?��s\.���GݷO�m��ݜ@�?7�A��M�E��X�'����WQ ��I&�z�8������xZK�B!�DmNg��ߜ�-q�.�&8"�,�>���HAU�u�`�� ���W�`y���C�#�e:{�� �-���1��D�[v�0�H���Z���ķ7�=���V½C�$A;D:*��oW�Pm� �fP��0�F^����D���_zX��C<�Ң칇���?���3�
a�yh��{^-��8/�Xa�!��bL�Aޅ��h��,���KV�HIE^��(�7�R�n�N�67�f@�'|������m�'�
wd�t�q�ǉe�.!���q�I�.�*��F�;�����Y���݂9ڛ�!��� ���'��(f�.ri���
��`|Tg�W�w�Й�M���6s�e�@(ӷ��=+y�g�
�؊L�Q|/.Yʐp�?ܙ��ԝ�۬/U]�5�:M���n%��jz�������KN##/~p��&�@�,F�bͻ
�jy?���=�|�O�^����>ծ�=d3��=v��Ux`^HI�R��`��°^]aJ�G���=�x���cq��e�ُ�[��{�)��^���g�8*�w��HbV�֚(rf0Z��±+ ���L%�H�0B���wj}�{c�Ңfo����G�GƜ[jt���E���؂��P6;,W
&�>�R2��ci�1ޑC�d�[�!��`X����l8��b��+��G5��8��1��U,��L%��Τ����������UiѨogR5�K��;�W�|�,�+��d�	Cuq����\���ִ(9���#p�;�i�	��]`o��F	Ya��n2+��a���%���uR.���<N�@�9�e�:
ʮ-�nZH�Rd~mL���I�|���GNR�iD6)�zG�~�h�'��.*5���ʺ+e�M�S����Y-�Ȕg��_�9�ٴ�2�9ϼ2
�;7�|Q�3�O��0��}��Zy��o*9ݺҠ���*İz�΃��a�7��t�R����8ԳG�ev��w�[|?4 F�|�Jr��9��g΅���h�[���f[�}F$ <�dU�ȯȂ���tXe������"���p �����v��MGn#ッ���Cq��Y�����P��V/
3[-)d�'k*��o@�m�3:؏��2������tXNlLg%s��826_�C���"dO���X�GwD����n�͟�:?���E��,f���J�c�珬�^�B�*��W^�_���t�5o�&@&E3��Ȣ����-��ؾF{NA��X�~*�óVi��N�m٢��p*��B*�$9�D��zq�d�h0	��Yu`b�/��o�k�s$��z�3͠? ��P��"��k��fTN���u�B	������ ǣoy�-���L���G��� ��\�TY��^G�xi�(Ŀ6�:��@�����d��}O�ν�w]�������*	�f^I�����v�l�ʑr^�^`���+�o/�V�3ξ5�3	� ��8�������FC��6�B%:�^�l�=���7���[k�?Ut#�5]�gC���|�䙘.�O�h��c��o�J��N����ݒ���֤یE1�sA~[|V6<�İp�k>��j�vN|���8��qy�rƘi����P�\�0�u:9Qg�����WS����9��Ɏ�k�S�4U�3����@WT��q���|��Ob3�p����,�GR����(�x�%�	>grO>Ts6���aM�껀(ױ���:-Fe���b�L�H�e�1��3v߿Y|`��$�(�I'���&s�ĩ�[`���?֑ݒm3]w�ٙ���E�w�<��\Un�ue�OGo�	�N�D�X��q�����&<���o)G�~��'I���8����U���c�|��Fh�k��>��������yOm�!3�K1�c��<Bvbb�*���n���=�P�³B��櫮^��8+�������pzն`��fp[!Y�;p��W�׹?沨�í�Q���.ނ����Ǥ*�V�!���O�x��)�55� �~&�਷����V���i�]10'vd\/zQ�"�[>��X;�	�g+fX�������ؾ��Q�I�yaYB�E[H�����De���K��bO�*�W,k�}j��r?�cx΂��S ����e�n��J�:߂c���@�Y=��9m���4���MX��^��)h���ي������4W/_�L��ۮ�D�D���T�^�$듲=�o0��|U�ɊDk�5�Ì�JL�~��
�C���jLa�l�1�\��S�&��1����h#���g������yi
t�jK�dh̝���A�p�uH�審*S���nt@�;�;�j9j�й��&Փ��Zi|pt��Qq�{��R�M`x�6�T5�1WZ� �[x�x���(�&z���~���K��চ�r?��I�[W|�`HϢ�u�QU^�����)��5t�*@��'Kəz�{3����I^v����c��x���?�7~ǰ�UD� �q#45�XS��'�UY��D�a>��J%>޽Ma�t���kY�F:�f�x�m����G� ��A��՞ҥ�ed�����Z�
y�AW(��1'=�yo¼?��A�&���yX�S8�o~7��w�9�һ�ph߂]�?�r�wm䧗��a��c5xv�i<?g����7�^������@I�|Ʀ����r��� ��{��j��#�}�I�p'n;5�=��U��'�z�)�8����!#yX�fը\��^r��L	?�Ό�n4Õ^��G_�^<��l� �*B{�e�,�,%(�Q��q�s�iu�5p�$�#Ͼ&�oS�NC+Ƿ��Q����N9�01�TxS�B���p�	iY���\s1� ��\ �!�	�q��]�u�T/�N�迲�{m�t��F�������r��&h�_--��mB	z��w�����\�s����r*%8�i�����C��wݺ@D��]����F�3�h�Fcf�@v�JV��JZKx�7�d��B��[�g$<����z
g�t�b��mc~^�u�M���,��xH(��HG���U�߇�Y�����}@���G�H҃���x3�3��*�C`��T�'!�v���)h?\��
k�F#qY�	/0wܸ�IL�L���;���J���,��A��5�PoS���sd�%���A�+]�$�>�a��� f.�K���(��z�`!1�)I(mI����!1���%�־��H>�ϸqw��׻�#��#H�d��~���f� ��/�),1ؑ�'$L���Ba���� g
Z2�� `�(@�mЫ���dI��S	3������b�8�1�����m���$$�|��y��>��T��Ɩg��)22�"��OuI�H���f�ւ/(g����: �����,�<�{�`��	�^fw�g̼��9�3��_pC_G�ꁝ�tK���T@��Z�b~��?�������up���ğ{���/�|���w1F42�� ��ڸ�O��D=�1��G�ˈ4=�f�]��H6�t�}ɐ��a+��㙵e*&�z#�z5%���7�q�)*����D��m�+ӿ:�v�i�_��GY�,��U��X�^�VzX]��:��j�^�j&NF��H�7�@�%P�4�*�J-�B�നQfc�+7��r��ٜ���>ڨC�Jjә���mk��l�J$Yad:��'����G�=¹ZK7E$�	�$7J\أ
������L,x��k9%�&c��>5��#������1�֓v�Yt�`ʓQ���Y��&>�N�����(3�2C�$���.BC$P�!��Iى�l� ���۩����d3�]ݒRT#ۚV�.2�΀�N�h�d��XF����U��t�C��?���9������(O�����aM��"f> G�M?�B	��.�<
/mJ��7hd+���Ҋ�~��?��
�������35�%��a�7�� tbM;��M����i{$�m�G'��]�]I"�cW���jx cي�;Ӷ"����9}3!B�Y�M��%`f�՛�ӁTb���[������ ���b�{s
�<S�I�-��8�}p@��k�5)�G�����E𜨣���X{�x�?�A�N�f�.e�Ae:�"V^����r�\����"ٵMՏ+��Vq�����˫l/d��]3���'k����
��(=�:^t���SN��E�P<�P7q��X��*B��*F(!{N==������ʁ���3�ӏخ� �9�r#��=\H�H��5�G�ۿ�3�]�u���������ވU��糯��u��c��gq�}�S��oōo+i:MT�p��z�\Y���Mn����#���@��S���!�m:�O�Vn;����=B�v<�����y��$X�MRj-K+�����
�l�d#M_N򃌨J�����x�V�T�5p �:�<y*���?�"�C�衄��L� ���Z��ߧ{cV9��{7��7�8��	��k�o"����
� B;|���\�	U��xyI���A-��r?/��Mq�fJ�wR��w���; ׾¸-��erh�[5�u��<L_i��P>,�R�kf��, ���`o���9�mjP� 3@�
'��F���ް@�=.ث*�晵��T�������
A���i���-�4��B� �q�����/2�FF��A<� U�����O���G|�`�RA��dX�d����8���t
b'm�8�hG��m��Q�)�8k���D.�݁����%0����p���.iJv�;۶����������G���{:��~�oI��8s�QgQ�PqX�PTM4�ђt����c���� �cZ�Ho&Z���P'G��r5��(W�ͳ���������t��z�����ڈr��3�4�.#���Q|������qJ�\�j�������.3Mӌy��6;M(�q@�[��{T�u�\s`�q�D�&�ÞDI�ࢺ6͈i���T@��	����3Oz@����'N�܇sv�m����H0�?Jk�i.��%�栳���Qg8��@�����ąW������g�\�!��{u ����KA�B�.�g�D<���-�.t'�X4=\b�%��C�ђ y���qb��k�S��\
��1�A����V
k��Vy)�7�t�
�N��*���m�MƘ��|���ǃ�bƠn��-\fdaq���Jy<-{+8�7�O���qn!�����r�}��|���%"���fG)˜��=���ob��YZ��7�9Xn�y-�X��͕�p:�*/+s���؞|���y�i[�� |��0���C���	K����f��V�-����bK�r�MD��z�l֖�w��L#BCx��v�;&�m�Hm�ҧ\S	/��I��z�x�/�6C�6����=���C5��Zk�y0}�ƭ ˳��{�n��͸�~R^ �Q�R~��V��y�Px3��qB��9��M�Kf-�dU���%7J-���z���i��d��f�^��+�uz�\��j�i�2�-e���-O
������ݛ�W-9�Rz�)��p�,�R����
�yt�-���P���?f���Ԁ.֚���BF�6P��b@�E��#��
� � >�_r�՞�f�@�G������X�G�fek�@ ���G�K؄�o����4��2�I��������	\��hQ��"Dk��Qa�O�[�����w�m��L�5�	+'��������+\�ķ��ƥ*���s�a.m8����V�}$���~�4���?�j���|t� �:�o�k�ˤ�K��a� �N�2��;��˃t��> .�}Gy!T��&M�ZϨ���c�*ڲye�#J��k"��Dt������#�MS	�_�goR�:���W+�j����H�u�@�at�3�7.����`e�����vO���ޭ-NR��$��:��`4K�8H:`�"�c_u%p�#����GL�~�Pq�͈j�S�Eo���N�UGٱ+z�]Ua9�3E��-78�5H�!S��h8��I���\b!-/�Pc��x�wˀa�T�h�ҭ�3�јb�����_�Y�ƫ�펾`X����tA*����2�W�Jg�5�2M��R����l������_��PF<ރ�$�k/��sk�j N
>�+f�U�Q�)�	��YG<��#a��4@�L[XzeDܧJ/8��w�O��	3Ю(������_9-V/�zX���'SG�l\(5X�BJ3Mc�*��0Q�B*zD�:E��������B�A�6*O��5{������%��\Y�,��3����ؠ]��غ|�zk�42���GBSK�p�0$�dh'�f;P��;��h�i�e�L��E����t"`�@|�/B��\R��D��Qm��җ��gx�j�����ٜV��x��}-k՞�ͺN����J����BJv:�t	�}���Z� `X�x(�#�{ۯN�g_��-�"�e�gM����N΃#&�o���J��p�j�^����(^2{����.��{���v�����N� Hk�5T��;7��$I��=9Ƕb6�~����Q�POb&�ț�<�P�&�rk0��yo����> )�eY���5��vM4�Ú�V��~�[(]���덙��o�q`����24֚�Lj�Bl���C�O0�"����E��+�q�
�z�4��S��VS��|+�?Qzm�]�G�ن����S��\�@��EPg���|{c��eE~�q��e�����M��R�F� ��oھ��27A�0����=䁏�)k-��\s�IY�ɷe�/��(o��I���?^9	Ga���qW��]bpv���ƍ������ZP)ƥ\�t�}�Fs�OA�9%h�lbzp��[����^ ��^��tC�R��~��3c�)q�dL�T��C~Y�p�Q���B	S�ѭJr2�����c�'�z��R�*�@����񱹨������~7{ s�V
�is��b����K�EB������1 �`	YRZrZ�F]�����q�!�4�P�AqT�����b�]z��~1T8?��X���O���>T'�R>���!��$�t�6��\��]O~�Ҽah�	�LS������u�Ѯ3^�vm6?�i=��^<����I�r9U��徹=��֮F0I�SD+�pdY��陭�(�_��]�T�P)�F����%���}�@w]�Cx��W�����鏻M\r
���p�h$7α*�!�8!�]�`���h��s=�����e�1˝�_�`/5��.�wCT_I��~L�9:%~��G���sI-�iiʃx�8c7$�@�VYzs-!(�𠊦W{��{bT�fU��["���r�O�+�������hm�R_ظ�x�1�^���z,�:�ܨH��疊SeA�)���,�jY��\$p��-���������EweV�թĘ?<j�RIyN��1��|�\j������C8�ɣ�n�c� eRE��� j#�������Ё����Ɖ�Z2Jpa�8)�MXtxm�S���>H��{�V7.L�=�ˆ>U~� ��+jU�;-֐j8=��o$l���4�3��q��e����8Ql�Z�h/������n��yn��a�q���F�!=!|?�w�ޤ�u�qO'�� /@���̱�,�{�������
7���isZ�r\��f���ꕹ��8_��ޛf��3����BAM�_:�pD���eφ��\��HZ-����9��4�������+4��u۫�+��<���<���J�w;��� ��I���/1+s����{��]�~� ������V%��7�WAvY\����C%
�z<?d;�[�㏍Nr}|:J����u8����o[xd۲�;�i#�juJ���xѕM����E�B�,}����
ŨIˇdy�v����ZP���Xz/����ߕǬ���">-�Q��2�4\�g����^�+ڄ;�p������k��_U�e��VU�i�����zC]�bB��R-�棆� ����ژ��N.�G�d?�V*K�n\Y����[��AM(����dH�(���_��9��Btk���@[�cf<�
���b(�0L|��W|��(�we�`�?� ���K%jr����lK�\��͚EnN'�5j�i���]�Гw��ה&�;Ţ���Y����<Y��̖�n��G�o���"�zZ�G�c��Y�\�d����׈��(a�@v��*뤗��	/ZvЇ�5a�7�'�T�k-�w��-I��P���зq �ƹ�XN����xr�k�)�̱�ȵ�i��E1�`������|�}�MD^��}�F�iM�H�OW�@Q��&�xs�c�������[�h�}�F�M����-Y��~�-z1�.�φ��$�wd-Q�
bU��6�)�2�y#P�+ɆzR[e��h �b�'2��ݝ۽al`�a,G��"���2Nr��!s/]_dIw�?c/����z�?���\��L��2���ќ��~R~r��S*�H�3!��8FbqNv#�mgSg!`J$�26 ��/b�qף��A�F���	��/�%M�U�cg,KM�^W(�'e�q3��O�(<�*��f��͆��] ��zsm��:�+��+��p�'���+� 	��RIH� �KJ4I4���n���L���!��K��S��x�17����˺F�y�en�������q��`Z��y1��7�>֠�u�YNFup%�hٱ��kė���$Zj:���IU ���ծͳj�Y����+�����;����GS��!��֫�󤈼 ��<�8��r}YK�.@�E�'���o�~�5;Á��~2h�4����G!x���-tLDb�3G�0ڲ�"�7�d����5�wF~^O;�3]���6a��_J�j��.B���!f��י�1:��_E]��<i=|h�G}���j��#z��á_�9��.�F��"sU�%�
R�;�Q���]���
y�5�?���vk�"������o��J��v�~����%/���������6���.�Jě���%뉊46He/l�^�Q��g�=��[A��"�$ L��Y;}�&���{;5$�\1}��#!�:%siC5e4�]�9�n�3�o��v�EH�!�"��*��ö�sL7F|0o^Ǹ"4Hǟ�O㰤 ����%)ϒ��O�?�$`]]K�o�`;(�n6�����`EQ��b?�kaJ͒����6��ID-���,a�N#W�.�����9L.�+����I_Oܪ�I��-�7��$R�P��$^���B��6�Eӿ������-M����`���oSH�;<�s%G�ө�3�3��P�o�'�e�n���e�BN#�)$�)�XM�������ņ���:0n�u��Z�d2o�W�A����w�J[Jj����|e5�%�T�(��׵�Y��y�>|���Zs���P�5KϸJ`����Ɂ?�(������2��#�?#�G�@In��?,b���̲�
LG��n)w��=$�r\еq�ҿ��;!Ը�-��h�%��m�}L���J6��%us��pj����7�莨��8���
�PT�V&Q�Og �X#�F�o{�w�l� ��A��#Z��P�=��� D�����k�{��[K>�0���6�g¸^/��O�'����b6ʕm�c4G'�3�HJ�T�a��Yo�bL��cjxʠ.�6���R���@a��M�ے�b�3^гP�1Uyg���-M_Wo��Y�=�woޙ*��?G�b6��'x��|���f�@���Υ�孁o���o��� �u2b9u5}h�#YxҸ�+ �)]6�U,t`�^VZ��P̲�}>��y�_Pk�l�BN��Cw,o!�����q �2�sW�a�U����� @~Zu���Y:M�"�><����DHݡ���,��Q�q�o�;H�GF����`o�vX|�bC��=0�M�@��k𾢽*���
���%�w��n��45�oAB�!�?]";�B�������w��(�3��>�]@��[ r�}{����%=�$�����=��+�*,���n6���<]Z��:z%Ci�eB�ͪ9�׉L�veD��.Po;����dƠ'4�� H1�߀p�z3�I0-i���a�#Le�w?uv:�)�e���`�?�*Ц�M~�|)T�yx]] �MƟ�y^�S���������!�j3I�$�c�#My��t��N�=��a{�6��8>v���;+��}��%��J�㏟��O����".�Ypl�otc�E�jS�WQ�8R��� 8D�h��_�Vh{@��]��|��|
�ʷř1]�=��2�x��4	pP��,FIc��)�ϖ\�x�W�?�vӘr/�3T�x=��"ڣĈ*����2 '�n���FG�걥�[�6�V�7ǫΜ��	�A^x��ue���*�!��8�Q8�t~�����?���gv�@�{��e�O?b��1j&�2\��4�>�^�9��g�(ؠ�7'v��۸�,��͝��!�"�i��e�6���-�9W�����ZN� Cte!
1� )4�^��O�2tk"���:�Q��T�*��1^ �Vjgo���2Ĳ��Sٿw$�D��DL��W��c�l9��b�9�OrR!����>�?�Θ4#�u@� t5If��?X$�i����DV�mT�����s�V�~j���
�$t��`�*�\����n"�de�%%&��L1k��(��]hC�&BsN���#��X|{[_�9�Y־Y�P{��dW'-�s!���^���*r���m����l%6�P"�Nc���P�p�L�1F���m�eҮۼ|�cP'��8v�tߜr1y�4�蔉�Y�#��vߥ'���tq�� 4^�(���p�<�%�.M~������u�E�!����y$������jE>�H���ٌ}+֛�2~$�dVǱ��)V9��t�S�0�S������b��:Q�T�%B�vw��]2f �g/om0fz%K��r��s!jK�Ex����{�WLM��ߍ�g�WK]4�
�d`���}�X���0�����=P!R��(�=� �;�H����,pp��T�3ڻF0ج��,'+;E�3o�ߗz`��� �K���Sce���|f^��_�z�(�[ܓ�����r�Z!�;)����4�AR�H(�D'wmc��>���z��9��<JgI��>[����W����V�W��VF�>B:��S��Ȳ�m4p��K���L�_���5��I�K��u�a�~ߚ:f"��[c�������dZA��Cy}�l��PT���](��UY �`����Wrn�4Ui��*�"	�H��j�Cg��%7�7�$�8��3P~)��7hRJ0�(��Ef�(��2�:b2�¸JH���,�4Kw扞'Ne�
���.E'����ѡH��(!F�Y�(r� �(绽�)�Ϯ��wYi����{7[j��ë*�����T�ފ�8����f
_ΡD>{���vA
����<����[w
���q\� �K7�"o�0���Ù���%�qw�FX$�,�5˒���$����onɷV��e(/�c�ן��)��2�Si`�y7.���E!9�R��A4�b�׷�����u�\M3���L�K˼�X�HA;;ZH!����H}. ��^~�H�Q��F3�C5�M���kM?��G/��}�e4}���Х��I�N���4,�'ؘ`<S�d� ^���<�^���P�Q~�Ɔ����Z�X�s�bP��W��lm�_/_U�7�FΉ���H�O	����)�� 3�XI�6�S/�Gꂔb#�
4�{x�8��P�h�����*��� .�=�w'��ǋ��Bo��yF�w5�%������ɮ){g���Oݭh�����:OK�-�7���ɻyn�T&�3��O��k�Z<а�%���Wݰ_���It��?d©�>��'��t�f�=cOEF��R3�R%��Jl���]gE!w�K	��pd��r�9���/b	H�H��Fd�V�����ͭ�\`�.ibB�(��L�[��]q� �a���&�ݵ|�� ��ұr��k�堉�i�Y���W�)K�+4
v+�.d�	N5_[��ДQ����6(�����ۦ�nmg�t0Άv�O��j0�v���N~��4feช�cm8~̧���Z���Q�W���N;��tb�����N���^��;�j��%�BV�q����A��o�Ѧ���;�};I�u�������n�a?s9e� ����*2���}�$�`���#���%D�&r�#r�YT\9����0�^���0�Xn�2IO�|��W�lWE��?�F�Đ�%s��ꥅ��x���L2qh��n}Ƅ�y�W�Qp������l'm�R�p�6�0�<?ز�5����xumC�b�FF���2F���6�صT��p_͔���Mj��c��"gn��XQ��>�O�}�C# Dv��S���=���o���zk�w�J�~���LM�,�u�?�`���mwz7�+W�zh �|�����������>�7d�y]Rty��9t_T�>�ģ�DD�Ag&,a،5M�]�����T�er�8�	wl^��(Հgl&?g�����o��Bp�xl.��@�J��ֈ�_�]mV!�{*�-*$n���9�:"�Z?�e��9�������oVX��5���wM���&I=�V&_��?�[�x1x�QO�pJ���(�u�`V3������곹�MmH�O|Jbx�ۙ}��&o��ۏ�D?�����1����>3X(�X�D��E4�smm�������"��29A^k;�I��\b�Y@���>��.����i��3�J��J[B��Oq{)�;��@���v�>�ǳ�H(~��m����Eg�0#:���s5C��<�D���-��u��l�W���Y��/�Q���:ݔ�"�]@��J��N�0���U������x��{�E=E��H�k9���n�2�|?,�����x����?���@F��{,�������18x�Qyb{���l�X<��PE� �x��b������"���^JL~�W�¾<-�8bl����,MVD��ꎬ�X��DI�x��Ҏ �v?����L�f�X�~	rz�}&���3���>"�%�ߘ���{f�5����ŀ��=������v���53��}��bfmT�</�x��T䔫��b^�-K꡴A1�k=v0�����pcY��?�Z*[f������t�ճg����ڇ�=������T��4��W��:�i�J�m�f������le�}�g�T
"����b��9
uz��3�Ԣl��EB*H�<_�J�W�{�T���	
6�����d�T���!�-2��RKvU�%�NN���� �����շ��������#����w�`�	a�������Yf�7)
o��X�	��gS��ӭ�o�X��f0��E�r�S�(�*�?����w=���Q_�ڮ]�iѧ�o %l�v���"�,U3a��+?۩��D�@����r.��`&��Ѭ�J����}���w<����ֶ K��Q�V�� _�=?� ������ൠtœ��K  "�7at��_�D|=��p>T2mr��	H����ՅB��(#E|g$���V6�m3�c���8zy4�h���ͤ��LQ�����؈ӳJ�jJ�~��?vtk#��c����0�e.Xɒ�m�~V�(�����s�G�T��݂y=j�w�͉k�P��B��*�t<X H�$}��J(�)�GH��U�������4h�}��N�cb=��j��׈�Y-p�.M���kV$C�|�-�T�M��Pg�"����F6�!ӗu������ny8�U��Kٓ�Rm����C���A�'�;Ș*X�Z�V�{@���^'�J�^Vc��E���o��A�fs�=����e��R�<�|�a�צC�������d/���ys�%/�� 1Ge��N
��Q܍%��Q��wz#/6o��w$2'KަG��ʷ02��E��Ϛ��E�̙9c�y��w9Xz��G������7�
��"�̝���ob ��#(0B�(v%a"�L�`�
8��w���47'�^�������-o|cɗc~g�J5����)�d�*�O@T�ʜ�24���S�Bw�J�n+}9�G�So��E�^���Q���,��)m��R��eѭ�dΙE:�̼�����th�F;.ʲ0%.L�1x���weƏ�-8B�|R������6nMT�?��椄/�9�w�^YEn���v)b�KdP0���`ӛ<��� ��T
^g�u!��(GXh'���
�v@w؞�SI�NFu�B�� �ԍ�:���ڟ�F�6�*ϧL	6*"Ѹ�׍�َ����O�K������p8���?ϐ��;����Ơxw�l]]����W���Q�n?`�'����]�Jw���r��W�~.E�Q-�K��щ�V��ʓ���(�@A�"X������'lc����1^��L-��g3~ׄ���Gq�R�u*������R�m��}||�a( ��G��nب9M���
2Bʸ9E�
x��ik���U�`	���ښ?�%6߄y�N8���A*��LZ���0�h\/_�����{�Y���VO*�̎�.��ᩙ��)�n��$�kV�;�tLN�x�����G�O#�^���1��"��|�-��9E��L��t����|�ގ�_u���y ��3�[�G�V�	��B�A�$�_��������Ľ�/ޥ�x�~�O?�ݻ ����R
H�U��)+_U�xl���n�h".�<M�4��C�+V�5�Ð�f(H��F���j�Xن���/J�R�4h1Fjr��0��/�B��?Yu��?}Q�[���:dqu���d�f&{`�=��uFj: ���@�;��X{��J��Vr��F^x���y�+,b=(n��ĕ>,�T>�i��
�X�{���Qf��ղk導̱�tw`��a�;Bπ�r�xFH����nQ�ו�Ft�OB"�O��.�geo��8.��bZ@9m���Ő��a�����"~^A�	��_L��ѳ��A;j}W�±�,@̸�������)y�@��,�aV[V�ȑ�
���B�OHž)�$��.�~;�'h{1 �	<}�KF; ���W�)�ǡ��h����K~.;D��O�o}Frv�l�Z�L�	��`8�,��?p*�<���~��� �!pG9����Z�1��I���q������cN#��гy0!TSv�)��O��;\�7�]�$>�G��	��!:�e��6p�\�x%CE)�d�k#�EU.Vg%�p�ͳ��+�a;�,��꘭ClۄCnH�A�p�+Dr��1o�p�K��{��x�@7�ߕ{^�KA:5"�a��a��O[q	���V������Q=n�j�\B�}踝��ۇD�?����5�4��כW1v�	;$v��R�����ɺOWfp
*oMA^���{ɽ��(��������s!�)p�����rKQ��=9�cN��+Ѻ�."��ԕ�K��fC��n\�HMd���n���U��W�Zɋ*��M�.������q.4l���id^�M6Q]�ظ �G��Y��+6n����/,	��8�aq%���T'\3��G}��Т�yb��n�\;Q�HiG��-:�Kk�B�Q#L\Kˈg~��>@�;�i�\� �y�s㏂+D~]�ZΪ�ɑݙB�&n�u���\HWm����xܞ3���Q}hG8f�¤BԆ4�� N�x��b�J!�ϔ$�+��7R�{lDRlGZE�G`<U~�pO8�*W8Ʒ>�O;�>H��hL��'�ܤ�d���Ty?�}C#�'�k�����,���9?�����Ñ���'���ȑ4/]��W����,��	b}֙=3"�=e!#GZ�8q �'�H��3~>��@_���4/��d�?�&ܝ�D�W���.�@��Q��%��70y~��9U|O��L��
�?���tǌ����@p�W֒lC�7M�n[�T0~���Rl�BYɰ�5I���SP8}wS� x�PT"(���f6Z�FNB�&�Eͱ�Pц���3�����p�.��	
#��`/n��Ͱ=�L�L!�;��(HD�w�}��Y(�,I�Y�̿&uĔ5Y�tP|ܐ2��'��nS�3~(�y����3̘���&�L�;�zCV�c�Z��ˋ��:@֤B�&���c�7���\���)Y'����Pf�����"��$T��"����g��R�Xg�&*�(�*��ET��h�^_ѐv)
!0E��Z���9~t�8&cGҙ�7��v��}���thLe@��!�Z\^����5W@7*���������\��cY����F��o#�k'ߡOU�*+�K�ia�o�]MA���25�TE�)����X9<�-�i�%9��U;V�'U.��
�о:�uX�Mt����J��$��ۦ����X�, #'�.:��{�9�;��A?`|�/����0�T��O%�}�3��N�X��x(�ͻ>��KV�������έF,��lE�
m��j��Sy���|_o��2"�=8��|�;6ܾ8�*�_�G?���v���%��b���E��j޲�'l_uN����s�6��|�M�|H�2N|vs�A�����C�e=�.3���)���~�d;�2�2���\�j�[h��z���Z���2�2�u��N|��{Sn�z������B�"B�-bW�u�,�y��6��WL�Lޖ$f��|����Uxi�@屭'/W9���b������c�?�7��]rɆ(��j����d51������L]6�0��\�9��t�`��#)�M��w���Pf� ��U��t|`$Q1y���i#�lHK@���]���}�2��{��m����o��B��PT��������D��AF)���kw�8y�Ӛyt�T�;ϬGf�~���'�ˡR��>Y�?X��8�i!��e����t���>��GJ���j��x����-�M���W���w�kg=g�%�'���	�{>l�K��B���n�X��l��{�����W!��d�Yp1�1r�xw(ʢ�.N������ń��珙L4'���=��f������Ƞ�$$���ؖ����$���'��Q�_"�.fok1DY�v�GE���!G�xE��_���7��c�#;�@��gP]'�U����X��5����Q�,��(���G�]q�a�`����?�� ��Erv�D�D��E�
oH@#�3�2��
b>�Rr�g��;
��	�'�Y���AF�m���K2~��	G�3T@���O�u����i����#Oq�fPЄ�ƚOc��/1պoz`�D<33U���	��n���D�gR��t�� 4�1�$�1�X�H{�-�j*�Q��$��>~¸����l��%�m��Z�*m�2xr̍��'�-o����n�ݸc�C]���]�G�6s�,tD�bݹ�H&wH��	��L�p��"/�K��L�s.�������ԢϏ-����8X�$Y3U�s,	�F�2���R�~�w���^�������0T��8�����"�Q�i��Q��4�TE%��]4�P���nS�ń����Ջ�>�Ʀ.?G�x�I���9�Yh�`�a���.A�9AeO�
���jW��O6#$opG�d��4M��t��������&_�{hO�f��9�uv2�?�Yڔ��q{�mn,c�����O�G6�JF���� �g*��ԟ���/�4���c�l��d��6/Vn�C��HEqn@s��T���M/9�E4 o��noz��7 ����G��_�]$*E9�����;���P�)[�ۮ����3�_vI��S�O��	1s����A�
��~�?*��swH�rN������9�,�@	�J֍/PJ"�{����|l��.@��2�Gw�!k�u��{�{_�Y�:�'EFr�~{!��`�<K-�jg)���v�x����[ ұCuN�(}��{���S�ΏKRJe���YR�c1���P@���D��&S�nǼ���'�%S�c��Z�H�L�ŕ�N<�:9LǕt/Ԗ��G��|���$�%��1�XP�+m�c�x�\H73������q].�6��DN*X8�<�ǴYrɄ�};�E%��H*ǒ�Wln��"A% �o�F���S�v��35읺�tsEi0��3&l��Ja���z���i�'D�3�&>~m���)���3M
��߫Uh7��򛛋6lJ>�/�������lp�tղ5�T����ѿ�r�ʦ�C��X���_��E���y�k[2o�y�j����4�q�(L�)~�0"�qyZwQ�0꯻'c8��Ip�<=�����#K!gX��
6B��ƭG/��9m)4G(����L�e�3d�I���O�QЧdîGr�k�C�9e*���e��B$�7�+.��ߊ�[*R�fkA�s�}a���~�K����IP�<��a?\�������D~h�v�s�̳�߃9A|��JQ�"tJ�k����	`�(4b��މ��r���m�>���U�gj�C8�MC8�48#��E|�}/�����Yp��Qcz����l������rf�H*	X�%��0L�Ӻ:u>�<�m��.��O?�c�`���~�˸��z��穈+p�kz?d�I�X�sx>�$A�(mX.Y��E=�A����5�[��爲:HWCJ(�w[@�_��%�8�a�<�b����\�}~�u>�X��u��a���	��-����Z�bo\k�|���+�;��xə?���ҭ7ڪ�Z{�[�}$N��{�H�+Sm�$���!�y6ƙV�"~�Gl�rȋ���)|��j�X����R�
��0&�O����m���q�㌯۝wY���`���뺷��i[�P#b��L��,�J������3��,9S��ݽ5عV(�O�n{�Ĳ������v��F�
����;f���*]�^f������������奇�k@���C�4&���������;��S_}'?���M�ݭ�gT�+J���h�8��������XI0t��^׉����t�U؇�����q����X�q�â	�<��sP�շ��/v��氄� ���~��p�a�)`��?vp�9Q"#����tF+�Z|ĩ_��	r������L�ǖ=̙�A��y���y٫I��6&��~����n�ݱ��>? �6X��i&\���)P�%�إB���(�a4>��m�猳5ɥ���H�^�	N���vNVk~G�!tXZ����ĥ�-a��*'�RI�1�<f��f��2��|����]����O�D�[�|����������t��#�e�j2+QÓ�G#	���Q��Q�&>^���y�z� [��Gci�_�W/6;]��<{��v�~�1UR����S�B!	.��z�����烓�u&K�NT�I�$AN�)H%w�����1��b�b��Q���w"C�I�W�WC}�=Z�����2|ҋ���T�l��B�P{���+	�|H�5~���/�~:�����r�Eb*��-�H��`�jK�	P��?�U?]��j�^�/����a���U�-�]'Z�_�y����9����z}��[�������H�WBD��}C%��H*u�/q�z1J��T.fcL;�ʛ�D�V	�hO����tG��������� ���,�%��|�T����Ŋqt�O�W�r�i/t1��ɵ9�]l��WȊC��B��)Q�Rf�_��۪ÆS늙���D�,���=�YܦN�wQ^�]�e;�)|wǋ^�
�ć�/D��2�L41�۾j�F���;��jhDn�Zt3AU���L~H����wND*�5��r�u���!j2x�#�.�sJ3�1���i>Z���K6,t2b:�Y��怆~ �"���Kؖ�w�}-|�f?�����U��`Zh~� �n��l�r�ni���M: ����YR/���vA��2����ܙ�,��8s����΢
�%f���櫏�l�oF�����p�Ӷ�� '�L��Ã��8��'96:9Б��7t�����A�jċ&�O�����}�0�FQ����@z���ue�04KH�$ ��?ͯ2���[#�Q�(셚X�%���;bh_��Ȟ!��k��XS�`x �t/�0�a��؁��I�.���0~�)p�P��T,vIreD��p�z%!Ҿ�9�n�n��
s�17�N�(x�P5�҅3{�b��A�'R�vD�5;����I��B�Z�v�K�h͎XR%]G�|^��|�;�G�
�p�6��<8�Xې*w���eU��Nq��&�6R����B3��4x<.!w�GrD�T��+�G���YC$�׆��l��R��B����"�p �-���g&P�-�U^%y����g$�x��+��!�	h�$�lK�5q|6c<��c���.�6�e��	L\�X&�C���t�x�[j��/e�/:�kM"i��>HQI�Z���p�dp�` �����	qeI�CX���"!��}�z�U�l��v��(݉U�ꝀO�^��0LX�s���x��{PVc���H�^'\'`M>�F���w�s�ȴQ��t�:[Z�ṵ�����,'i���� lX߶��Ľp�*�X�M{NcB8Ei�x6����Y�G�c8��/�{��2J�_E����*53Cf�*��9�Z�u�8�:e�,�6R[�יFKvV���)y��>��nfRlhW^�d��\?Ա~�r�oc7�����}%N3�f,�!��!<��Jg�MhG`�� �T��1z��v*��y��b���+�-�F�0�ρ����'�}��9q�9�s}���%�8%��� &�o�N�%m_~��v{g=�Rw����^����^������� ?�Y��}��;V��������S����j�Hx�i�3X�L5�n���kO{ \K3]�1Z�k��mF�i �70��vP�m��0>���xn��u����:s�����L�N�����T��
�τW:��犛\��N�Ӗ��˗ӓ�֞��Y��k"ӗ�z�X4us���G �i�+�].�S������) ��':�s��k\_\=�=_�U6V�e�ɣ�l͔�K�K�0f�άAW�t�#�%�C��1{4�	�wo|9��@-M���KYɲ��s@>Km����zj	N�$��.W�'KF>ju��O�>�����ZB��
�ޱķ �;�͛�|�S�X��>�3pQ5�.S��㋡,1�%�B_�O�9�EOD8]{�|�b$���eUzN:���7���6��e%�e	C�	�����]T�lnW�{�T5�g�LU��ԑD��̚J~F:�#s`L����3�Dn}�o����׬�W��byX%?q������� �2������&���m�O�@�6�I�k�K��<��7�LE�ۥ�6�VN|5�W�k�i���0���źۼ����:6�:���R�u���I�����g�t�]���l$��ނ�3�r�+ `���3���YKC3l�$� ���Cm=��:W�.��"�
�8�0�),��Xd�4��!gԤI3����JÏ������j���\�����-�4��&�d6L܎"`��������湯z�K�?Q�e�����H��4C0�U�g�SY��󮢋bT��_dG��1���%�`#{�R���pYǎ��TC	���*�;K��3V-a�eB�EW���E��O���M�L�����,nO��kM�qD����S�B�N�q�)`�?�.Ie�d�[�	�B�̧0+�D>�GZ��ĺ.����������IT�
N���m����?�A��Rc�D��XwCC��t���hK�hwGل�zʯj�o@Y�(��@�EsEl��_�Xc��$�,A����{fmw^U΍_F�lӂ�,�%������OŌ�������Y[+7
\��q��j�����_.��Fiρ�l?J����y�a����NWN�`
!H���?��&��_��ɐ�,u��MP�r��o��O��r�[��]���3m��m�U*ʙ��np�~&iZ/h� �Z�"[`��5}}`b���B���]w���|�m��_���԰����)?:�0�=�gB6N;F�׀�]R�J�`�'y:�����I@�b�H�.'��2��4#�R���ٺ���87�U)�l��]�x#7�7I�׺��0�
N�Jf`(vɃm~���&�a�U�PgѾA���
ηu޹�f��`�8��jk�B���������(�0�P1f�؃��M��y��=�90�*�%��=��O�^>>�@�|R84v��N�pɷ=m�O��asTl�U�Q�eAa�Re�0!��q�<=��B|#hZT��]'�c,�Z,����=} ��.Qr]�HtH]�6���j!�p�֔�p������ȝ���|�n���N=	/�:�m^?_�b���P2�T�$�� �g�,k���+����P^� ��~�1�E�>X	H��:4��bk�z2sX��l���h� <��xbl�-��,�v��t�ܲ'�2��O��ϡ��τO�&��Op�bRz�~Z(O��5���س6�L|���RI|���UUv1�k�b]�j%�H�v���}�y-��_��ҥ�@?�m�oƸ�'n�L�8��4�abZ�s��U�=�Ė�c4�H"����E����8}���}֪5Z��4�/�T�*p+Oq��HtK��W.��& 9J��� �bH-!��̜GG�q#@��Y@!�4.+ d�s�3N��:���}��>בop^Nl�1�$|�_�:��vs�����T���<�]�ӍH��:��P��r��:<�lO���&����"����[���"Ɏ�¥V�P�^ﰿZ������Y��w��U�~W��Wdr��0sYG�~�^�6KS�lf�F[�KC)\�&eu��������U�+o�s'x��if��ݧ
�35G^��`���"MU��[X���胶�s�\���2o��HNA��BOV�!��XՌ��C�Q�@Q�	��;�R}w�D'f%W} l�D��K��uP�Ԝ�m�'v�J6�̿�Yp�z_���� ����@T��
�y i%Ԡ�w�ۀZ]*6�w
?j<�XˡA�u/N�և����VژT*�f>�4�z?�)���i#Y����xdp�n��7�|�$���	Ɥ]a|[�$i��}^�彘�����c8�������i�焮��h���B�BJ�hYJ����^��aƾ�i��Y�����fYIn1{k�uR*^���p��M3N����Q���'�1�w9�Z�~V�W�����o�=y=#���"y�R	T�O�D  �����W��>@�e�E�� ��c��R�d�H=T�$�>��'n8m��[�;rc���#�i��
��3�0D��㸯3��<E����q�<y9f�,5{B�fg~��*IL�=/|��B�PƎфj�0���[������`F9�.��&h��&�,��F���$w\JB��O��6&�y�R�JK�0�f�#4/�`��{׾O�q�w|��ި`AP��]\6\����r�=Q[�S�IR�4�$�����s���z$��ڌT�b~�z���1����`��c�wAIde���#��� n��HUfY��N���94�Ś%�.=z���_g��L�"�����O ��Y̽�S͹��i ���I;�l�9�4���Y�9��5�/ެ�0	�^$���������*�N� ���_����A�]L� kw�c�R#+��� �0�"��#,8����+\h �*auY�����s|�%+?[�ʝT��m���(��R�͑S!^�]���ᨣ��^ҠL�Ѹc��wGBf��_YS��}`��j���&��0>�jY3���}��M��1a�_����\	#�u;G.�b�*TG���[i�H)����Y��&��C��MY��T=� �
�^f��5���^R�sU2@R+!п��	�,�g��l?��=��I�1W}�[+��K��==�Y��+����|��
;�X:�K��l�rE>��P�D��LGS���]���������~�|�ּۚV��n��!8����N:���{lX���k�(����q�"���G(�q�Sy���Q�(O�/A��c)56���V*���t^�'�p�z*��p�c�f0�,{�|�Ǭ�e�b��-6�|wL��)���;�*|9��󽄬�iߒ���S�����Ö��a��dk�n細ڗo-�U�H]7�n�L+2��T��x�B쌐N	ޅ�K�ׁmgu�C�-�B��74ԓ�K��Ph�Z% �
����r1���VȨ.	.����[&*�owO<
��ccc@��2�xB|Z�@�����I�G~m��v�GZ��S�����~�+)Y ��-u�ܭ�k���_2�t��[��Ng}�(�$2�
0�:����s�Mb��y�����Ȭ�m�����Gof���!����	��/E�4��'���F=�\%1K�����6�pׅ����D�F�Q7��K������J�$�82��.t�b�Z�B�v�x�&�qH�	݃�s�Z'��vF)¿Mk)��]s�dX���FVeI,c�:��<��F����	��I`!«V���zĸi l�Ƴ�U�e�C�}�i�e�M�e����j�r���4`�'��#�ݧ��_��!��*׿��ߋ#����Z���_fD	�L��ЖB�f9�ǵ7�&��12%��,�n5<�|���G�gx�� F����,_9�)7s�e��=L����X��*7׵X�E�8$ȓ�KF{ě��lE<%2r��N�ܧK�0w��w���T^-���38t�]u�"J���
X��hiB<�]��|��E>6a0m}f>?a��a�R�fcnd 4aK�^~0b��]�R���w�.�\��0ou�V9�I����C���.�{�10&~e^aj�5���7�Ȕ�g�@DZW&5�{��='�$3���~&PcR'c1C���(Ka�����؟�XL��2�K06͙��������W!���p�%��rҌ?�;���c��7=�����k�����J��w��Pe|mme�8��~�x�	�����*��υ���{vOi�Xf��Z� Ě����K�>{�7R�T7c�q^�>��r��a�����g�bL��I��gT_E�d�_=��rO��.��{�*��?��n^�V
w���n�"'�}��T����i,��������:��I���Nt0
��W�<LyM�U>���%�7F�����.}<���K@_i�AG�-|_�P,ϸ�����8��M�F��@)�H??��QE20]�o�����$�|��J�B��ƛ��R��	� �|0AR���_�����J�	d(�#�"�j��j?�z���Х�}TT\�����-�ު�x�ڈ����y|ۃ_�j�e���1��@I���>�f�g+0�c�I�A�A��R[���}g1��۴�;��.�������N�	�{c���*�����@�*�3D��ZX"¸,�Yf1�I\fM<W�2�y����[+�
�>b����Y�XE�yCy�(�-Ϋ~@��9�~�F( .%�`+WB'�1�e�_�N(��\�[H5w2�f<[l]�����&?g쳄��ƚA���Tv�fau��� 574�j���>*� j�a���L���*��3�86�)z�j���35�z�o��)��m����j�f�5�+O�muHk��|n�˰Rup��2	-#�K�㉸�:8S�C�������u"���-l�?qf-"�3l�3�0}PB�<mɋ��qO�:K� ��&j�T�)�=}����؄���lQ��H�=����;�&���+G��z�}���.�����++�m-s�B��Gȟ��вZe���M�oP��1eJ'z$���!� ,�|�\���׈>K������n4U�BEe�����jJ	\����5��x0�%�fJ�m'xy���ѿ�p�=����R�0����W	�x��)��4C�C��w�dn�DV?�&T�zA��Ψ<B��Yv�� c>�d�g�9g��b�����N0�຿/�1���hwG�4�lt�1��i��|���J�./�����1E��7��a	�f������ �ѓp��B��ڡ��ن��#��AF�l2���ڹ���F��Z~Id��7�I�lV����[A׊��-�yVg}4%�����ՀQ�G��t7jAF]0x��T���y-a~�7�;Dp��I�:��2J���ש�	��ca��/Ҩ���P��+l�ic*z�80X7q��p��hŬ����Y�$r�aA�u��ֻ����Ln�ϗ�
��7�\`���4hfQE�X��es$�V�����c$��heǎ�J����L�Ʒ=ii�Z10��K,?�@��L�$�q
�$?��21D���Hn6��mOB��'٢)�S�i�k�
0�`r�P�����!m.��JN�FZ��2��{Ӑԙa���W<�EȠ��8��v�:��	��`��.Xy�(�&���45%krp� �m��C=8�S����t��
/�;�|y�y�if��T;����f�oϏ�˺��cنt�f� Z�I�<�z8�^���5~���s-<'Z-�o�x�vo�f��T����P$x��R�8�ywd-*FE|��Ҡ7�c���X>��������>Aڠ���DA�}�u$+I�v��[`˂NjU=�&�Ԙftx�O��W�V/�OK��צ�,S^G=dBg��z�����D�ì���f�^`%,1N���Z�Ly��t"�rಿ� �|�}+���q���"��3��,�G�k6`M�d����<դ�8�C�-��f���Qo{�b�� ��u��CCk}MO=�.���O��
���ȸ�A���/e�=��-�Oa����$a�����t�H�s��)���F&�O��x	�$O��gvb������V���Z��1�����၂����I�׭ݚU���l$�����8��
�!�z�9�3y�f`nni#��ǆ9I�W��-y��r�t���Ѭ�����ɡ�m�������@��1r~H�kV�����C�ʯ��;Mhƅq�?���iP��K��͍�W
A	&��f�Z��^��'��N����=5��@����G�ew r�F��������>k�?�sREf���`��7���bl��Wj�ua,R��>[ʪS�Kl5(�b*��~�
4�ǒ��}ՠYUd����wA���x/�k,��A�?5�H�3���v-�e�BX�꟦ڮ��/F3�9�u�a�N��6uR��O���5�ȷ���L�Y��䣅�����N��Ł�:�T����iLTܪ? *�2FV���Y0��LC���B�{���u��齽���u�v���ZP�T���G�gʝ��m�9	cJ�~؋�L�B�����p�#�L,�	`�� 5�6�p�����}��&���1*\����Eґ��M(O{�}Tz�/�ͤ"�v�ꚙ�M=B�T%���=N�`�%U.B��c6ǂ�6U�(x��R�B�'��_ �C��mZ�ɓ�(���'v��G�_�@7!��>-3�������P?��9�v @g�c�-��ŋ�G'WL���#�n؜��I��PT.,��qhh_.,K#jPػa�����7��ug8��c��3�`��6��s�vظ,�<W<x�/�*lP�=���tQ�,��6�4�<�@`{=Ѓ]�c��I���߶�@1U��oξK����L+W���ތ}�&����w�23��\�8vE}d]�*G�@�A���tTH�9��OS���ֲ�nE`�MHLj�׻>Ñ ����՛x���X��1��ͽ��Cw�G;]x'eT�E:'�;���	<�<�+�Ʌ�4X�ϔb@��N��eaz�%C����]{�er���S�R�,�N� ���	>N�2S��QQoJ���Ǡ���+�B©����豰y	t�~��3��#����.X�b<<��_�̖�A��N��2�(�,��E���B�����Q���ec��[b.�v�N�%G��%/�c�����9��Tv�*�h_M[����˂�N,|-�1���d4����E(.ˑ	�
[��ߏK���^Rf��=l�PQ
pc��������C��U���8~�<�֩,&�/&���v�Ӑ���uin�t��k���nǚ��X�&B>�ΐCY��"���FGbx���(�it?k{���E�ք�VY&�5ν�Ny�2�����ڤ�q���V���]$� ��#��-Q���؏l}�
�yb.0���Iq��Z񨆆v_* HX������F|RH��E�p�y�t�O��V��o<c�6��`3#��\��:��ۜ �X�����u��:*�W	�����'/<D5��ER�c��x%��]�c�"�ɜn3ozBզ��5�lW�&�F��v��!��q���2��%)30'Y^���V��?6����,���V��%����І����T����U�������Q�}8g�~��������#������t0��8q��`�s~G��F؋��
���Ie?�g^��_B3�f�HG�@c�z������cI	���5�W6���)�����N�Qd����Np��#Et����#�\_�ǽ���:�� �'�}x��^�.��gb�V�g@��MXۣ���/�ٕE�Ƌ����T�N��o5�u9-�o!P0Ux�cR�p�����|�^)��(�έ�� �Oz]>���`S���Քl����V&5�)7��_���l��ȩ9������F��y��G����Rw�{C?����ԙxI�:y�n�>C�Y.��Da���.��z+�W�t���x�4�*�<$��)��+OT%^<RH)!)�ċ'J�tG��ߙx��s�*�m_�h)�v��;��+���~6���`���v� )��������������8��rR�u�Ԅ]C�CO����8�P�'h]C<b�PS�V�N���ħ�&��UJ%ғ�4O	����c�����m��i�}*���!֍n�qm��xP�^�;yQ'~�l	!Rݾy+�C��O&�ڻ	��Z�K��@`&�2��\�1s�؛`�NF���:���7��$���N�nQ�����8 �ek���1`�6��.�J��tb05����G�t�p�h�v�/�%�ŽRVS�
>�����	�$���ӛ���5h@r�y�x�} }?*Wt�p6��Q�&�0�Ǉ܋�9�{�*z{+�rm��.��tC*����I:�&jQ�
��ʢW�<������t�~E���!Kr�/]&7�#˶o��fڤP�εv��N�L��Śc\d���/�@�X��i.���K����4���f��������.��װO;����K��jy�<(����Uώ�G�x�%���Px���7���^��xἭ���!0�8%����k.��-�v����i�G��<���m u� �4�C�e(g��+8/�7�npU)�A;��.[�>�Xr��ұȢ&:�-�yD��5k�)����G���������1[n�NF�bـ��N�{����b���ѴӁ��6K�Z�_�����mU���@8>�M�e@�~�w2�x�"}���e���x53��^�O�v=�:U=� ��l (-?Ik�"��8:�p=� �[}��$J?+���J�W�ζ>K\F�}�������N�S*��E?Q:�Cd3�B@�x��w=�,�"?s�yn��F��bX�BW�3��g�
~V���^~|c���iB��u$_�M:�Zt��Ƃ
��]��O��b^�I��-�����`'(���4�x	��� �ͦ��E�?�&0'�S�غ^W�<�`������~�-@��k[��:gX�,���/݅
+���Ľ�rK�w�N0-����j�yB ���;���������#]N>0`�m�T�lh�`$ʕ������B��=b!ԋ/F~�l�YG.BQz�$�`I���o%um�w��`�f�w�A��@n|#%B'�hpF&s���1�>R�&y
e�]�xO4Wts�ҥW�`��x4�^�Ij�`C�c�ʄ��������b�%A?HW�R:8�+h==I>k�mk�0
}���_B��p�ݼm��Z���pB2�D���
i���o��O1��;g;ݮ���4?�\Ǝ��]E�볥����'�nr���הrxR�O�͎�0O�� �������a��;b2�b�6j�!�]�Z�wP�y���c��n�G�G���4�{A|�2�<�Ȩ!M�~[��:;�s��*��8�Q�(Ӆhʞ������O(ǧ\j��z1C&=�6=���٦MS�ȹ
�	7\���^����Y%̠ƳS�}@������	����h=�m��p)�������A�uWS��u����g�e�m��2AB���T\���t�5��׶�6�d<�r�r>��������@��̪ɀ�z�{�GJ,��r� i�l�~�Y�?���^��vw#���=�����K1k�Dv���;�c;��f'���u�����{��Q(������ ȋ�w�V4��_�z��6�ٞr )�6��*��r�7[4g�62m.Ɨ���	�6���C��"��&���zÎ��c8�����R��`aߒ���\�#�UT���,��T��d&)7�0�-a�Ǧ��,����1c:����t�^f5�P�����w��lCSj�I�o �L�}JiB<(�[Y�s=��ȯ�q5ȼ��_ίf�˱:c!D�'4�r�<� \f�<?$��p����A�Ƕ5��7�B���NXP�˰1֎ϱ�b*�%B<
��](�i-|OH�$�b�g���������)�P�i���A6`�ő�ǈ7�sJ�b6���rF���1u��.aZ��P�E(�1�w"���;B�-]:���Z�Mv��#�G��P*�q���LI�aH��~]��h�iÛ��)����	���16t�>o�|� ��8R5q:��V��A�z�0�iRZ�)���)pq��?~m�b��'�;��}����Vy9����L�o��������`7�6�i�Z� ��c�Q�	:؛�R\_�vk���߂���$tw��)�X������!�/�h�SyfU�'� ]���\�,,_�K��?R�m�6VN��MoLl;�>�����(���M��$X%��?���󹇳�>����~�Ǧ��� or�q\�N�m�7Dh~;���G�����~¢|���q�����ƛ�=��I#���:Ny�߉ɤ�L� (�"�1�K
C���}aYi8x%er�T�p�t/}�	��r�Y@0����Ew�n*7a;i��T��w�#/|��ښ\v����ä���.�T9k��]���3�`0Y�[�����44N�-4�%�⛰����9}�q<��r+�·q;��Q�.�"���%��[�e��R�Rŭ�����]2k����!���C��*i�øR�G��I�}�Tq,6�4���F|Jپ���
��C�Q@im4��0�$\�%�$���g �����S5WYk7b���z�bwb��pM��Aʃ�>Պ��������N�Ϯl��yˮK��#�Y��e���'ʛ��@��E���Nc�)�	� ;׶�=�{�ߝ�jA�&��@.�+伬�b�v���\#�]\��d�c��[���ynȣ�A0�i���-�炱9ټ��"'5��u��I�C�0-�Q�l���J_�;�L����b�����]&��Ib?��p˜��%G拀xkx�9������3�aѡxS�vu�d[[Z�3��?�
�6�5�j�o��U��������~��vK02��"�FG�$خ�Fâ�3Q�H"`�f�v�<�S ;�:�H��;�9%hO�^�m碙���DGM@͸c�V��0,��NQ�7h��q~HC�d�֬.�P�EJL*�W�=��B�8������� _���*9@Vɜ�8=�zr��`Þ��7	$���9o��0�z�,H|(;�'�	�P����E y�\�D�X�a��g�,a-��a���L�%�0����+\_�7��ACltQ�D��_hV����k�\xe�'�gF�rB��j]4��z��#ɜH��rz��3?�\�p�>��M[�s�O���Ars��܈sf�X)Ռ"����L,z)-�,F���q�ٔS_��ż�X�;�J��:%�~���7U��)����@Y�м�"�N5����7��|�z;�jJ��%�d�)��<� %������ ��	��^X���ӗ�fǧN�zAR�K��(1�)Mԫ:�W"W��vF$�̠�b���9f�b��~��+D�X}o{[��B|7���.*~�v��������7A�6��)����S$pO�N�
�|x,7��rx �=��.�T��O���sL�8�Yd���J��Қ��ۀ���:�9���`t��UG$�>+�u"���4s�7�~����itɪ�ԧ�7��!*�&6��y����y��E�Td���8\�Z�Ι\����7ꢤ�LA�Q\� �Q�AK�պ �z�t���k����b�\�:1�voD�����Z���V�p�{���2a�N��7��ٟI<��}݃I��c�"���r�,��)�"�Ͻձܙ������e���ڡz�g���.�t�s��S�׫J=VF���C�;eGR�*����V�s�W	hҝ=��S�0���i>�͔�I������e���@���x���%�bZ�<N�m�|�0q��5i����t��3� m.L�Sל�r��8��b�&��򺍐|�(.'���qx'�{�}��>��e
�Y��2�&��W,F�n��F6�*�¢<:�j|":b���J-_�R�cc�_&��!T�$�g��BےPM�Sd�YYA�ѺAa8��z0uʸ�/��Tـħك�=���)�}�Kշ���f�]}wk4;�� �/���������=��JA��W�Ѽ/�[�W�	�ً<���#��.��d�{�H7!��e������������\NߘN���N���]�5�|w4n�ݖ&�W����{Wdٖ��L�`#:��VB��d�ly�W:�Ժ �}�DW�F\~�	�y��L'�$�Ƚ-8i��D�Y>.
}�2�+� �rz�FF��h+a�ۚ�����xV��D8E�A�|L4g���U���O-l/�`&�
j^�'V��1�xqXw��Ŏ�m��t���޵�����,AH���*��|��e�.x�Z����y��y*~F���1�\�L�x%R���o�����Gަ`ɕ����*��#S�����ČE��1�GLg��H�wF�To�i6�9Ӿ�I�J}C��d��%����W\*w'@&Ú���70Y�Y���T���ٵ��&)�S���л���o���`���I�n/�Y��@m5 ��c���t*��lo���%@'���5��#6qa�2(�^O)q1܌��ޟc��a1�e���ݐLa�)��%e�5fPJ<t��#�+]���i�4�x���s���lN��㼷��?,-	HU�C]��SH��=��.�Z���df0!�I��R^�r��ԩ��k�����L��91@�;�F�^BЁ��y�RK�|��+D�ӂa�!
�59x����|,���ۃp�+�ELJ�q`��	�o͘
⎘���mWU� � ]X���\�5l��0���߰��8��D_]=��_�g�+� ��&8���JZ�`&M��o��h,7])���U���/{UԦ�tH;a��#�>7�,t:�o����%��[�3�S(��&�"5���-���3�YOVÏ)*I��It"����������(W�UY��hP�:�y�RWgW���WJ�f��[��cv������R�d�Br�V
�����6�-:��3u����G���ud��4�Z�P�$�����M�� Z flW>���5�]��JW�ٯ�E\ ��C y������U�b*~�vg�n�W��̹������.%vm>�3��x����x_^��]I�wϾ�s>�@��z0�����{G���T���'`�í:�v#�u��rV�B�CM��g�ؾ�h+��y�e6X��t��\�(�񭵡�GP̗�hM|G����-��~��]�qEr�?�/����֍�A�O��+?��]f.��w	��2��vF�IK`"g��a�SV!�2�\�zW��6�P
52�3��k鱲�$�M��J�p�r�qP(Ꮱd���o�:])�N�V��&�yyHՉ7��@�>�|��ǹvv��30P�(5���!���Q���`��6�c��o�)�Mvlj�#*4q���Z�fΞVڐ�!'Q�'	S��e4]��%R���u�J�� U!Z�"TUȭ�~��!�7ui �{p
e�T�w�R")P��}"���g�tX��V$l����`�;ј���%;�O��Iެ/!]�Vs�}.r���\H{Y;��PGlG��E�j�xG�ahY��1�����!�3��q� �Ĺ���/R�9*�rTFSM��6��B��mB$�+	w�(��pm�FZx��A��|����ׄ�g`�P����N<Z��a@�U ��>7�+t��`[��@$d����E]���Lc�4�K�AdT�Ь� <�Ve��f�ϧ\��O��(@`��n�_ �{�d���a�lM�5+���"zX�<*J�1`J���6��T�Ґ�
.�^��!D�,0����>՗w�bw�kY�X\ZM� G����$��)��L��K�J���ˏ����pś��P�0�<@�0��J����~���-�-K����:�F���#)g���)��k;��HąTs)QWk�}Y;��T7AYzܝԯd�8�����zD�����1�_�+2����?�}7;U��~�	Fh��t����5t[�oi�������4��+�y�2bz?��"�I�����4�m9�
�����~�<n�t]b��J�~y��m�X���7`������eD�ˈb��d�}:�z�Z_�v�g�P�K1��~[�������H��a���-����D���@�R>�*k{p(8��c&ܒ���8|dѺm
P���Ξ6�z]�F�-iG'ײ�����%�f�T���U'IG&0�ZT�QO�k��?O���F��-��$���H�6�)�Qv|q褗�Y�[��x�A����9u>��6c�l�b��������7X���Y���G��C��f����`o�,x��Q�� vHh�W���}D��B3�PV<T�~�1�R���'�
��òhO�T�{xʔ%�Z���X.�����,'.b��9��Q���1ΈL4������K#�$�2���X8d3l<��zǂ3�J��6��i�KJ��z��'mn��(snlr��'&y�����O�t}��f^�O�5�S����SZ����򁮋�a�nUZ@��%���2J���Ʀd��p_*@ɿ�^�öV�+���1���C�F��³���d�@�sbQ|U�SaJ�Uj3�:��I}@��u��Xݵ��U\΢p	�w	��۷�[�5:��̧<� t9!Iv7�~7�QB��oǨ�Ǯ1�R�;l��X� �<}|��/��{�n�&iF3��AR��"�O2��Rt׊S-�������/Z�a9���Xi�?�E�'�'�Yk�4�L�#�8ID\u;׆č<���聵��F)D
I������ջ����WJ-��Vٹ�,i��O~"�+���gxX��2bp���

f�P�� .�cґS�4��XA)G9g����� ٔSo�R�r�~�=h��,�{�9L����FE������٩=�L2K��A��*�g���/X-�VҞeJB׆TD��[
X9�2�$��V���t>���%���_ks1*S�4�Bβ�7�LBt?{0q�4�9>ˠ����?"��m��-��6<|?���z�z7V�a[��� �!֨��E^�	9)0e{E�HFa�&p<}a��@�.(|\��y��<��Z�NTf�ǖ�I�C2��!�췯��O\�&Ӕz�kO���[�[{����Ν2\�F2Q��A,�yH(�jI0
���>��;jQ��"�X7 ��q�����mF��a- ��E!P,�n����-��{'����u��p 6L�,����M�-�W�Hdx�N�F�)�5�	}ۄ@�6�2CvE�U*k���Y����ݾ�u4��,���=��ծi�B��rC�����%�����v,�YT�Ǖ������E�8�1�.Aɦ�l @$lW�{���'�+�V��[D�*;���Hj����)���*Q`�H�lۧ��>e(�UP�ǘ�"r�9��{��3��W���?x.)F�d�0�)�Z�.)�{s�	��_t8v s��^6�z ��-9������V_q��N3���ґ�57��Gm�/5���LG�o?`I �ֈӷ%Ѫ�
�M����p� ��0�x��X%��BEucN��\��z@��~�D>k��N�3���]�!����:ռ�d�������c�k�Qo�Q���1-6�_/�%���/m�_�� ���۽�*'��F�]#́0��ugۯV��Q��Օgw��z�S���2��v�C삆�Sm̇��_�] ~�,�Vȕ0�m?-,v�9��|�(o�
�<o���m[��5%s��ҘB��:���-<���Z���{fT�Pj�[�����G%c�]���� P��o�]�5����c�s1����_'0Pꑄ�R���������5J��g������{j�^&A`����
��b��|�,M���;���=�)Aq"r1��4r��*��5/x�������.��!+P�O��"?[�S�2g�)n�����OK�K�x� 63��VQ�_���bC�����1c��z��,m]l%@�M�q�#$"0TO�uܼ��An�t^(����}u룆"�G��D=���l��&}���g5mrOcc;N#b+NW�3�-������Y�B�X�G'�~�s�`!Yx�PfR��?,҄Y�%�>÷��+��B�}�����>ٷ`uW�dk/��T<�I��Ί�ʉ�(�#h�H�Y�y{D�yX?�WF��SP�lR�xkK�)�Q�M:�(��.x}w�����L8��P�?y�8[�s���:d���f���!I���[�/4�u��?	��A��Pg�������� :0&�a���J�q��������`�O5�4����5Kw��ʝ���.U�˿Q>�j1�i��tҔ-M��� ��z�*d�9)R�G�_͇g������IMy�ϒ�w�}�G��x����⺮��%��x���c����z4)���|��.�x6���&cH�e͑�P�d�T�� ,�:|��<��W[^�{)��&�Q��y~��q  �|�����W��	#dB��!�v9k{)�hY�{��;�f}��=�4�l�غ�c
7�)��Q��\-*������8��]�<�4����x_7��A,�9~���P;5J��at�\�ԧ�Ⱓ<s8n�|�*��Q�{l��k��fVڶ���ĶQ����� .h�Py8�*���7ȹ�E����/U$�� *�t!W��J9�{�\4�f���P���1ȰN36��Z�)�\�z�0ħ(ge�/��:���FfcE"_�E%o��z+�N��.4��t3q[t��Ȼ��~1@k�<+�7:��0ѹ%�7����"y�u#6�FM_�p��7<Zq7".�f��4;�]�Y/>6H���<���\6TQ������P`�L�F~���Dڻ6Oc�5�:FA*3�����M;�q�fӔ�����P��7-�*�D���a<#���ۢBb�U`3�+ExIzd�s��#	��N[�����Ӡ���'�:\��)�%�,����J�@�\q��z��nV/K�y�l(z�D���l������I�jy*�P��|ԇ<�7���s x5�U*�5�k�>@�^��%fj=-�%Ӿ��Gy���EG�>���y�mzKW���*�X��1$��*�v��o�6�H���ӂ\�,f�Q�+Q88p���M�1At�o��hIxcV����E>�]�� ��룵����������!ތj�v�zkm#U��_]65`r�n�<����<cyJj��HH�4���Un[�V_�;�DL��K+�>�wc��������V�=��cW �Qe�7��� u/P{+@�d�=��.�B�X-�� �������Bc9�����"*�bd��
U!C��E<]�F,�!�v��@����v{���&m�}~�>e�D�^6�z�H�t�P��#�8�v&�5	<W�%:Xl@R������U���˨�5WF�hd���P2�'+�*dk��"Ne)ԪeI��0Mn�
J��D !�y� q������zhZ��M2�v�Y�w�gv�Q<���o�q�!7eF����Wa�Ɩ�C�h� ��p���:�ﶾ�S�h�����nV[L�bW|w'����,��s���r���)�V�CjU�q���x�P�PM���(Ð��mH4�~O���|)c�^kW�vǖ�}L�$�!��b��EZ�g�x���5���)���A�$�q�Ή%�� ������;z�s����e�q��}_��M��J"BLO'��Nf|Z݈!u��H>K.	����2�N6
2h�Y�z/4���j�/�B� U���h��Ð8��$#xx��Y9��b�L�1��2+iV�i�a2'W���x++����� s?�\�uhG�;��Eƒ�
��U��a�+ נּqtZN%z1ˢ���"o�g���bi+R�;��pW�OZW��Sv�W��2 Ոl�ɾ9nrƌ����U(D�����P����j,sT��/�r�۟h�S�N��'5!�2��	g��藎R�n��2�U�R���ʯɷ�r�� ��PW"7��O�t�vy�FO�q��Z>D�;�O^�<t�Y�܅n�	�+7։�|��A�7�
��k��2}J����h2ԁ۪y��i�F 3�Da�-���❙���Z��#����Z=�3���R�L�f�xE<-���)�C+��޿��y����{]��+�j���ď��pŌt(�ۜSG,��
Õ����p�QZ�WaEQ�7�#~[�����R�mRQ������Tc���L";��mԻQ�	��񺁟�sH�	�~Ǻ�B�3��Wvy��R�̏���2^崤���:�D�ۨ��!�򬗧+���+����:g�d�u+�n��ʠ�^N�I���&���c<��#v�=��e�������Dh�_���Ku#���)- S�������BtE���(fA���]q���a��`]�*��o����#ulw����b)p�G��������-|�pp�d[_����:aի���0G.�1��`^^�����FWw��/Ƹ�@G��:�!m�E|��g�B�P۠��+�kg�O��� �(4-y�l�ݱ�u��S);��z�']U(I�,����Y.�I��:̦^�gG�+g��6�㼺	^b���֙�Q�7����?���H��h�
��e�~�XK��{U����0�èhUzO�m�}�]�l:bL(�2��D�g���vӉQ�?ۦ�u��r�2�^�7�[���(�X��7�
���/F�2C�W��҃F�ä�����T���S����{!�z@�:��Sl�o�_�� ���X�}V��ΣGH8�\������)H�񮑘D�ˎ��Z���=�|�[�&��� ުӱ&�K�*ZNb��� ��X8\y�[�*��斶�|�����q�>��"����p��3�)��sO���b�����վ��\ӑX�H����[;[��y��6��g�sW��gE�c�^��A�Z%6葔��
hv�����֡�d*�G<��oDb��f�"]�5Z��y
0�0���=��5�����3�$~b�N@;�y.A�C�D�_��_���k.�5i�,u�Qz���ް���#�b h�5d|r	��n��䠪�~+�Gdl�ڒU���4 ����.R��ꋩ�]`sW3�V�3��N	�j��Tl�V�P����1�-z�	}q.���;lO���S�G-����(��Sb��%�\�t '����o���-ͧ\��	ӕ��F���a#>��=+��u3!�d��L��*���K��^`Ɖ���c��7�č�G��`w�tE��nH#C�Rv�n|Ǣ�
c$P�����azΤg^�2�0�s��_���z^MP�s�̊Ǵ���B��ySX$/q�C�!���s�7�>���S��U�@o���:U�>Y4�m��	o���|�|o������P�̝ѷ��X��'��u1a���ᬝt[U���ҥ�H��1��18��7��+ʜ{��D%E�������n8^���gNG��Q�I��G~ ��N�{��{��*��p%�H9�S�&�4����f��(g�ޮ/�&}��.|��?�q���'@v��UY%���n/�@Q�
�&Io�A���"��t�@�׸puY�&f���|l2�n����]&����va���L��Ήy���Fb~�	-��!�`����2�?xR4P=\G|��oQ�sV�<�RVu�IZ�W��@�Ml�A�og_x�t��ֳ{rnD����Uw��bd����5eE�L��c��Q/�Y���t��#f,�Ya��K�q�t��ݮy�+P>�a�%|�rp�����3m�(!}��o�:H_轨�Y���b�>f��Ly����s�ߣ����L�,vmaTX�7:�h�K�M��'4Qeʜ]WGo��S1���k��t����K�튤h�h�J�����S� �]R9��ۺ�O����ӫ�ո�����(�Ls�+��)E�ꡒ&�e�S����I���9��(wq �m�\�LE�Q�h��|�����>�ҕ@�B�Ԗ����(��uCF�#/�8��`�UJ��jM<��}���|O�{l�te��4!�v6M��y�c����?�<�:�]�(oZ�����;����|��Av�� [E���'/��Mf[�u��8�����-���9�Pg9�N��''N�p�}KXY�xbh��햓��R7��T����0,���|b +Y���� C�%{?���Q���Z�T����B|�F��6�F,v7X)�ڰ]�d<
����Է�]�YH�yo+��减C/+"��xȅ��`*�6��ݷa�)�(#ƷT�bW/a�z��+��n�B0R�C�R��yyb��r0�.!��d�F�P�4s�vtUO�+�Y�L�F=���Yq�7���ߞCkoh��3���4F0w��A����&���12�ڨ�K����F<�?��(�,xg
�\>=���Gnp���ҟ�g��\d$��5�[���nCۈti��"U�R�j��%���*C�I�?��߼�xH�X8��ԉ�8V��#�����I�~y�֩��a�`�S�,)�Rm�g��8�9Zh�yT�"���F�\�^S�kS9*t�q#�"��d�N�u�U�N�5]&��3lY��}F82?�K}\�)�2Fє���x���p��jӞ�
@,�ۂ4S+���m�6�@��ڧmzB�7FN�y�`�Ľ�~0�N������og�<���\����@����6�x�o�B���i�n�By��!�	O�rS�[��$��vچӑ�թ����;��s��$j���LtC5��:�.1bGU�?OQNOd� �(��x�z�^�S�J]�;H��攍���L�I�ֵ��!|B{j^���ɾ��ic���P����)�1;���i �|���W�LF�B/Se7d
�?�N�\��mp0�0���*~�}JL���GJ��P:�RF"<Ew��	���zn��1?�j9����2-�8Ǧ쿒w��$T���T(�j�S�<Uژ_Wr�GV����NN@i��
�,�a�⮲���7G�co����/�j��1=�x������ge]��ӷ��@��y?\����~�r$��9�bih��k 6�Bs0�����I��?A�<���+�Qa�i����^|��+�W ����T�a�(�_ۇ��
�(3����c�i?���}	�g<�e&�i���6��;���yQcN8z��-��[>�� ް�yQb��0��@(��ݰ%zْzkYލ:�n�BM8i��G�l:�d-b/��?
&&��\ϭ���t�"��(�7g���B�QK`T�{�V��ۨL�0\�b�Ę� u��F�#f{L+��m���l,!�Q#M��c?��3\�-ê�lm(��+뵆4����r]�%�׏e��B�-����nv�����3����6��T��3U)��W��i�A�	�oCR"ל��8ѰZ��|6Crc"�Y���(~�d��͔�4��&Rt.Ǘ��@qP�ZK�~ X���w����I��HQr]+�Ly�N���ϗ�nt眣t���dSGS����6f�Z�0�U���z���6�'�������_ΐ ����W�|P����U 5�x�֣�^��������66�{��m��Q���<����Om,�r)�Q�Y���I���d��^<�1��o��I}�7�W>��Tx�QJ�F�#�7��䍢p�R���G�]��T�=������\�`d�q�Q>�'��Z���u5O�Ջ/�|
H��"C�-���B��M�.�ݡ��!h�	p�ǟ}���B\����p�6���ʚ��n_�fyMp�����%֚r��mb"r�I{�ok	K �D5���#!�R&�զT�C�U�ɂ����ߴ��l*��j���/
�po��|�YY�������e��i�;�`�ǟg�5K
名�؄�7�-;\ӆ��l�3~�Ԃ �dp�/��tQ����մ��z�D�ˤ�y�+�4��IJ;T���۩�[����j�����ū3mcN��x�t!r�.���8x'�aA��uƢ^����)���g���i�̞ ���Ś�?oG5 ����2�BL�|N��'?
�6�&sӷ���0�	B�r�R����V��an�)e0x�ƚ����|,F�(X�ϒ������u"U�f}fn���8����'�!r��.�X�E��E:�V}�	�| )�s�
g�������-�1���M�@^Қ̻ �~*�8�v��{�5�J�V�`���sݏ�t'Kki�X�E�7 �7�2(=F$m�,ؤ|:�K!�ʶ+ڡL0E��{f�f����)Ii����D�*\��O��>J4.ǺH�nT�v�=^2�J�)��d�s�Z)�m4�E�t����s��01����t_Y��>�������b.Ӧ�K�io8;�#�&���ԝ�>���\y��$��59m����>��Y�9J��,E��0�0A?�|?���}�X�N(e���@�j!��O:�<?�4XJ_#�3|����w��������	���~��B��0�~��E��U�6���G��w�VP�pE����Ѳ�9� �R�Y��P��n���`�㴥�p������{�B�]��T���7ʪ�<Dk'+�Q�^��Ǳ:9�=}F=�F)�_�@�9�cXi�D�%K��ö�w���]�.z���~F8n��U\k���VI5�'�]�=�_|�9��o�q4ᕶ4��O�PmQ<wM��
ʐL!>���#w\r��(����K��B9�����@�`�V�!���"�珲e��uo�B�1��qp)�ߩ���O��@�+`�zHV:�-�h��ZcBDs�2�ә&H1��xC��$>+^�*g�H?6�Ŗ��;J=����5%���fo�P��[{����O	E�nAK��y�")��XW٨����$3��e�"� E�g�\�S8*(t'�ˡ�8QpR��l��5O%#DQ��n@�əR}���gh�E�m8����xTf�Ӽ�A��=sM�Z�*��Fe���l���Ё��E��4'2��[�0��H�������L=��1P7e�]�-]n��0�J�_B�S�j8�4;#V	�~�=��}a�7IVT�8pNM���X)hys�Cb�/$���)e'�u�S)]ٍ���0�Q��Q�Fz��Z�5���Q���n�E�`+2Sc�����de���Ո�Y�����c�N��;)W*���)�٠��س$c�,xlG��_p�^W��სh`�T�_�zq�%M�bÿ���R!*`M�f������d�k�oMW���z���J�6�.�ep�����2����A�ފ�lh�!�G��te���g�mߜD{���<L���o�r�=F�%r9�]��l2퇊��Y=�u�ɒ$*���4:����쵭���A��G��s��C�\4?B_��b=Q����S���{�T�9�Z�ҥY~�:*O��z�7�ڼ�b����e�KM�����1����|�6Ҙ�e���\�k�j���n����t*j�7��7��),�3����Neo=��%�/��(c�b� |�r����vBu.Rw���7��lVh'п뫞�ڑ+
��`}��jaa�C�Mn�
0�X{$г<oז>��ܔ�d��ð��]�k�J��@��Ed?�M�u�l�NOr�"��1��L�2R�r���00v��L>8Q���L���*�0Qt�������Az�,9pawSm����ђ�����+P�*�y�����|MTJ�S���g���пƻ�3}cӟ�B�{bu�~S�\�f�4v��������rb�c�@�������R>\~��������E�ʪ?���%�#G�}�NP�w�A]`.:e��`Եt	Db&�R5���d��׷�x�zZ�/��Y�L������v4ށ�Z|b6�0c8��
�����z��|�m;��s���=�]�b��A
 n��4M�����Al-]�r��K\=�ͯd��6uK"m��/���O��BQs�?/��>����C�7=�U�>�?9�r���8�� KNx�]��-U��V��7�?�vv��N�MT�S�#H�p�w�Y�:�蜡����&�L��K�9�06)����r�������3�&�ykK����a��w��"Y�@M�w��	�J���TJ�����Ǐ~-��ǵI�1�ыRcnTm��(�&�\7|�Ss"��S�e�VQ�F<�ۏ��Vc��P��l.�>�,"]�I������9&	Y^*5�,�4v[(��	�Hw�)l���+mg���2�o�����ȑ��*g��d�ıs3a�)�r9��i)�L�+k��C��Jd�f�6N+�6�+?n^ݢոW��F5��ۂO0G�6w��/�x���m�oDbNsPoJ�!C��ꆕϱs�E��(�?��Q�9}s#m���"M���WX
���숗f�y�0đ���T̓���dg�IM�|�f�J
� ��Dz9XR=��PQNM9eB�[��d��~��`ųy�����쏾��RZ��5S1�pj O�z���y,�����Sy�yu��Hp^�}�Wí7Cx�cn82 wX�5ehQ�;��������L+{Ǹ�09�-B���*����j���!*�'`gvJ����+����3I$-8��)s�X�6�o
�Ƶ����3�q��@L#�� D��1���j��z#Lu��F8݁{r�֬�Kew.c_[��W�Q��Dg��6�Q�4����l��kz�**G�i����$����U�S�-��Py����'�d�9�ؘX_
�Y���@;������t���#�����FڧU���͋l¹!��"�K*k�ŧ9�_|���6��B1�;;�d3��(����m�����}Q�7 ��~�TR+ȋ�%�ti�%�9���SN��J�5# ��HEe˭���"̉[�xc>{ܶƏa�� ����꽱2���@1|��iQ����::���KMxc���	��ʵ�'�u?�G|��W� 8#��~����Sg�T�����=%�:Uyi��.��z����GZ�b�P�Κ�2�N#_�g���Ԗ�F��C�c�F�0�"�:[ֈ
L�`�2,��5o��E��8�j�b�jqd�b�{��po'E�%�`�\cu��5��� :�e�� ��>�~l為�]�����w��C��ͼ�*�+���[�E�Ɵg�L�ֶ�t)u�	M�����n��#7Z����gQ�̾ş�pH�W�;�����0�����&�8���#ـV�	Z�(��q2��d�y�=!akL��!e�d��%��R����ƞ�jxs��xM3��0ƕl���LW��#nQq{�f������(�{�b^C���wJ�r� y�>�qA���}�F&1cJU֊\Ne����8@���y�g�wO�z@o�/�|�Yv�$�x���4��+Q:s�z1�����T�s4j�gG���Ȭ�JBW��u��@(&�k�����s�fv`�5��c奥�mQ1e2�S��$�홲m����<8*K�颲*��N���� 0�������V�WHS,F�B)5�j���Q\��8ne�;lN:�K�O*���鷒��ּ�K����$?~�A�U-�"��
|�^���Y���y����߰&����'��)�$�.�|�����/��V�'���6�V� Ŗeט�{�������i�g�b�L�d�gC\E�T���W�B�g��<�`���)���j8ϒ��򴃫?�n�����x*8I�A�|�A��.o6�?­�q�҆Ș�Fʼʿ?�M�Nո^�e�G��6�l_U[��E��4&�����^4N8�W/5C� M�/2�O8��:���Pb�Sǳ��Lҕ���!�' M�����Vr�K��;
�r��"����a��c_�ke��8���Gx�81)_��ߖT���˩J(9���0 �3�	�3Op�1Gd�{'ܫE䋩���S����h��_��L���g{'�.��j���r�&Ϙ�Z]Ɯ�s�w�k�c^5�+��Q��P�T��Q$���>��6��LR�m-oA��AzJZ�|5W�Ҷ#6)��YF�6�5�6�ܧ����ן|y(R�\�s�R_JR��cʨݽ�����;Ǐa%�E���0|T�_]��$�1q�fx)49�AD��(��T��%'�2�=c��K�}�B+���C5���Dn�2K�n�$����8��Jk��O�&#ɜ�j�=M�����hC;6��|^�(�ֺ���@F�e�K�Ѽ�]N\��x����w�2�})xO�d�����~����ܩ�4F����!��䌖/tU�a�Ѥ��8]v�$�_�����D��T9�S����OLh�H'�V��j)�ڬ���t�� J���o��`�rc��|K�v ��.yd�H���������?�7�+cT}��[����G��S�o����� Z ���7�DJr���0lVߓ|e�T�?K��w���e�@��B@��
�W�}��5/�0�_"�y1>��1���o�m�J�5�b#��3�u9z����fb|�!+y0��Z> ��w|�[n���l�씳$�M���EMx��n�~�@&W�C*�x�0�_�!�/�KE̕u/n)t�,�/oT�����έ�'k9�)B�0���p���̔�.Zk~0���)�m�<HF���?q~�;&�rDB�=���	�,�AY0�0�Ԍ'��u	\����I�g��ɷ�b¾�A�M�$�}��	[O ��xXȯ3�QC��
�J̚�:�ۀ��Uv�Y���֜ ���7Ei�4�aE2e6��ې{ҍ
[��7�:��at�"�ɵ�ٯ���ZP�f�[)���V%�C��qڵao(L����a��{�&9�C0�g�6aaK�)'�f����C+�6L.ykoh�ėכ}?��G�(��[��Aw�_\`�jJ��YJag%�H����[o�H�F����@��Yo�r\��aξ�N� ��@vb9���j�#j����_�7ŠΜ���e��%8�b�����{(���+��s0:G,g���S���|Zˉ���~�!BV��Էas��\�:��� I�$a���t��QȚ2�,�T�����de��^zx?=�媸ף��S��¡air�&p���\�W#|G�	�I�*H8Q>�D�x5��GQ�<�W�/��D���:����6�k��{,*�b[^s.$�,�I����n� ]Bh�e�y ���)N�Jr~8�D\����p�ԉ.m��Y��㪉�s<��R7�"8ob�Ķ8�'So!BA]��/@Q�:�A�*���o��Z��֙��X���������U �RH�U���Z[������u³�v٧1r�(���6�*h0�ؗ�:R[E��[ˏA�����| M|�(�LRl��a(n�Z��hg1 �}RD�nn;_Az�@�`;�=oKS�NϾ��5���`�����뎾�c.��C��vN�_�|���^(!��v^�E��@p6��1\|j�f�9�\�"
�+	݅T<(0��I�24_��w���]�$�I՞�+ְ�����j{�b�נi�͜U��ޢ��LE/��Ŷa,R! �m�;�����K��.�[��‟��M2�"�	J�+�ͥT��Fib��S&��"e�mW�_j�_!��m���t�&*��Z��.h:��o�I�����^�-�������,`���XԶW�N3��,g���+���Ŭ�2��m��E��x�U'�*�0��
/�5�i��`�h�II��i�01���O�lgnȐף,����>��^�1���W�R���[A�t�nr�����Q�I'��GMv0�Y�1?L�~�3��Q@`�M�=? 1����C:��	tOKy}g�tD��Շ�y	X���������ū�`;�!\/M��,��8h?]V?�a�(2����O�y#ͧKN|V�	�>�\��%�ͬ5�w�@�8�H�(&��PR���D�W]�:)L�Ӻ��C!j�J�c�=n��L\��c�^S,0�rׯd�p�a�.�4�-m�0���~́ě��̙|��g�ʉ�D中�W�����7Zie���(�z����-W0�sY��(u=�<�'rc��8�ޑ	�ʅ�c]�����#��B�W1�r�`��\S���U��$U��O|�#d6/��;��_��ߘ���*�����FPcԲE��ŏ� �n�+��U�3Z�ƙ�[���MX &S�r�I��j�-��k����QjEO�>3n�JNWZƩY�i�JP}��G�ȝ{z���}9%�p���
v#�S.bD��ֵ���ڄ~��T�$N!4>�����n��D(0�sV9�y<S"�=IiX!c��P�����6dXW�K�Y��ۡ��s���Q�=�"�Q2��/\O��<	��4�o 
 ��:�EM��kNw,��πK����G� ��,��@����ۡ������F�G6�zg⭦+q1p�K��$FO�>A�ΰ��sEOi�L���=�+>�;Z��u{�/W�a�+��u{h
j@��T)�����c�px��p'��E������Xn/����U�>����/�z "'0��|ER�G�oA�5\yi�v�ՙI�"�2��%f��5�M��H}������V��ᚬ������]��C�#I�+M)��xݡxR�+��KU��x���b��Y�^��n�O�Z���ښ�Ս���T�C���t��&�l����#L9����1�=�/�x�qW3=LڸĪ�	v���Hc2��!���S�r ��аH�z'���+K�ﾩ{�b��?�¨�5Rj��D�]K�����@�#�t:ǫ�3A������z�+.ѵɩK�H����ok.ɩ�|�ڨ	7��k��aF�R�y.<�Q _p\K���H~x�c�D�m$aI���� ���C�}��4Ni�j�9�G���䗻:}��4]�+Jn�����S7x �Ok�`'��>e��6+�����$�z�a��F&�g'�h��� ��f���y(�F�k���Gfʢ�����/ݫd��h����/�nah���+a�]��{�������ZY�WeuK�s���Ċ2�ĮF��{*t��eV�ⰬM���A�Pf�����L�1��4�u�o�f8p�Y?jL�~��%�%������s��;�a����%,���xWQ}�� �����b�Z@� �ړa�2�
:��j#� ������ {�J�[�T�ڽxl�.B��%���,qт�f����\X��0���Y����瞹g�У�ׅ�OXm�5-"�w������!���}����E�@��i�G6|�\����h�.���J�)y%�4��W�h�H+h#\Y�FZjzj=��U�M�����%nv��Ѱkh��l�NM'�s͊�ad�3�G(�v�ϲkƌ�	���gŀeF���L=��+sʿ�w!�`�ea��'�TV���:��S�<v�5@�8����Y��GUT�Z=c/WՆ�uɟ|t@�Z�x��ND3w%_�"O�s'���d.�Q����������p-�]�R����;P��}�;<�>(ahedF���3mN��h=�V�I�+��Ct|5!H#fx��#�>߮)���h�뢖Cn}#
�b����W�r��n�	��6�V��1W�n�Tp����
g�LY��A�l9�����`��p29��[�s���m�v���z�\F�h/I>�/p��_�=M�d쀆l�RH=$�'yQ\"dv�HAږ�c)�l�>b�̪�;g?S���"]���n\~�B��G������
��y���.ns��C����G)�ՖA�R[�'��0�di(&��2⭅�C2���V}Le��{�ۻ.���zh6���O��^��':ڽ���8�HUD�z�0�X��y<jK-��S�ҏ�[)�v5Fb��;��S%�̽��*%��˻�sFnT&{ⱟ��X\�,�t{�D� 2�]a)��:��Y���u���]��6�Y�m���,c��`]��o�h� �����n���ؤ� �����1Q�@�K�	���s=��*���^V|�sA�wQ�ɜ����p�02]<�G��=	9/�C�}�z��᳆,
�/�e�@���"�f��Q��2\[I���7V�t��c_m2?Db��H���!��c�����S$ �Cָ�MXӿ~�����%�N$u;Ɲ�v�v�{%la���˞�,'PH�U��d�ww�s�(����A�yWzI�4L{*��&S+����Ng�Hu���jh������<(3w�{!�U��+L]^�<:�׹��ӧu�!�YWc�6�Ǖ�9{�ώ�x��D��
 I��e��8�d~�*��v:>��(�P��@MMϬ��,�Sj� �i���$F'a��}l��b�6��jΫ'�$Ď���6��AN��
1�7.O�j�(��]meO��|Qxw{�uNS|LT:�US��szO��� �/N��;Ώ��RIۖc$uB)����":��#�I��? H�9!��0��)��_����⭹�D�ڗ���\�8�E�4�Sl\-����[�t*7c�b��4����õ�S�s��p��� fb�u>�=	�V$��IL�X�(�%f��	a; �܅�	V�[R��I[.���u��R���G�� V��A�.��D(a�Z�!lhmozJ9)ȇB�3b����q�N�jt+,Y��--����-���U�D%�4�,uV��_`h >�ϰ$�"lگǙ�Ǜ�0F-MgJ�����͝�z�����?�k��br&R(~>._�7��^�t(�@sM?�Ykl)�Oީ?l9.������iB{ܹC_x&�a�����a-��Z4�s֑f?<��;��w� �����&5�b�\��tno�DtirW1N壂U�E�ʥ�b.Q�ߟ���bjo�n������'�Y�ђf��\x��ș�č��x�{c�!��.-Lt�c!��j�z��"��)�i�3�}ɸ�K�}R�� ߯�Q0E�5 �k��<�������~��H�b��l��U�sX����a
��D^��ӇLkD-Cm�X`��4~&��N@9%u�H7_�-6�s%-�o����!k96�>@.$ݥ��J��Np��s�-��Y]�Y����[Ar2�27��* |7��c^�Y{O��V>���$���w�jO*�a`y�~>�@�������H 3|�M�[M��6۴6�J�}�椶?$rњ��>��ӌy.���3vyKL�hJ;�{ӛ�+�f\a�$���Ҹ1"Wһ�'SJz(
��%�JE�zK�F�I��!i��<�S]	+��;?1��:��Lli��- �tgkpJ�h��ל���Nݔ9���ϔ���cw���15�������˶��m	��4��Ns�.�2�B˦DR	C���Z�s[1E����M�<Q��i��|�B��p`����X�뇣�|�E�.�����˶���*�]���ܻ]_J��M`�����?̕ξ~�|�6�����,"L�t\
&U��50�\�� �=s��^Ue��,�4�b�7��1�U�s��z��������@�e>�l����:/�k�����qX|I���lN^�-�R��Bj�}	�CC�����n��Z��O^�/�LY����ߵh���X����U�̌9��jψ�Q-w��c��̶p@�+��ř�9B[u�Fa�n ����d佉�ڶMeG�L�#��)a�� �W�XD)�f!2��*ߪӥn��G�<�}�y�L8��G!x�e ���=
�3m��c�=JJ��Vq-R���M����u^X?'���i�H�Ɔ��C��_�bkN��o�Q��x���@K�Z���$2�Y7�͞�e��W�-�e���X.�.��u%�>��x0��%�B�r��_u�Y�#F�g]\��-Ox8�@"Ξݢ2.t#�S�v�T�I�3ܚ�i,]1�A��̗a��k�k�����
�k�D�"P��ܶ������a��J���q�Rt?�"W�m��"A�1I�.j4B	���Ĺ����1��2Q��e�� A��&�9w���#�|r!��I��D P����"��E�pN���e�Ҝ��`[�ZNU�@��e���
����P�Rc��#��hW�y�����3�*����<�%��Ѯ�{�il{x�:]��L!uݒ�MI�l�����aAb%
�2Z��# '`B$X�Qa��b*pu��֊��N�0k��t���`��hV/�R�ݜ˺�"3o���;g�۬9�B����	�]�V8���������@%QW<9����$e���6������6�V4���G�5!�#%��%#�e�j�^��vݖ�U�TL^���E�r�s�5K׿��AuwU' ������t #.6H���G�~4����|�b�5��Q���EՇ�X�Y��lp�W�h���V�I�8�)߳�D�3�[��|�u��gW	N%Z1SJr��5q,�~�.��k�1J@g�h���	ʼV�Η RU�$��Z���<�+L'�Z�b���R9ż�G�� ��V
A���."�)��E�yQ��|���e$|�t��T_�4�tjj���J�M��~u~�%@�w$�����Mb�l�u��3U[���:��������q�_��}s��8;g$�؊����bC�#�F6;��ė��ǶO��~Uy��4�ҺY�ww��'����a~)���}���֥���s1�6�0p��TB�,�9�0h΅_����aXD�ħɵ��M����[���vd�Q����b6�(�M��i�T���$IP�Q��|�U��D��`�F�ϲ�2�8��P\����U`uN�P���˯�ec-4�E�/]"�^x<����\���X$�Ǟ�]�k��bn����6~��驫�@�4\W@���
"�D��Ԟ��:�`dY�e�ݟ�̢��$��tzB��r��Q4U`�r����M P���2h[=a�mώ�~�7e�������3�������O&?t�u}/�`H�yu� Ω|E�hB<$�6t"l\�7B@��+?�ڭ�Y*@#!���ح��15!8G�0ZnQ,���$���s��1��t�@�{�p���9P�V�	P���l�*�R��@;:X�t��E�g4�tE_|�'Ǽ	��"Ai���C��>>�
�d�_�w��h,E���+��7M'��D�TEG��h��s�Q�้p��?`75a �݄[`�A�øuχ ��m�����%@�c�5�UI=�CŖ3+�
�a��sy�]�ҥ:����v%yF�-7_�_b��+�[�� �١���x��m���y?y�D���:X1]�^Ĕ�M�X��{=��]}2;!�2��j7�<�G��թ���C�"2�u+��t�we.t���kg��t.�4N�`_�pi�{�94>�:%V��o誢q� ,�[m6j�²ޱ�P|E�S����)R�}�)���᝕fo�]��㞇`��h[���w�1�o��0�+�Es��@k�O��4V�h��Il��I<�
N}�g� - nZV��b{L꾔gT�(�V�?�����'��q}�S'�s꼂@�|�N�tnO �ٗ�R��B
���"S�eDi4��~<h]H��;�V�2�ݔ6���(
��092���0� �.w��cYi�Ie�8zS�^f�>�FG�zJ~"1�Qۚ��a$榍��S~�>^��=3�G��x��\Wd`N�(f
�t��)�l�]��𿧕�����Ɩg�ۙwCQ�$� �v�RM�/�2Lw�
=���t{�x�٩�W�.-gշ�$�
n�小R��@���+z��%	�)h�{^A���(�� �7�/���g�<$��m��|^`�*��p�U��06�9M��ߎ���s|Y,%!���΋�S�����}g����%���R��ا*Ʃ=�6i���9�A[u�e��Ln!�s<�?j*�Z�M�L
�R�)��74�˾�lr�}A�żX�������V}E,�߇=9�f��@l���<�_��N��h��-�f
�O$��EG>�	z�-��:�+?n������A�EuN��#b}�)����H6=��;(I��ٿ���{·=��.\R��k�_,*��)��b*߷�Á�;�́\�L]���X���$��Vr�C��D�����In8]�/"�-�b���b�C���ԬG	{T$�6����=�3���:7S��uީ������q�4�+rAS=*��eZ
4�'��j�)�1������|=�# ���x����������@	W@o��^`ŖgŲ;�dѰ���X�M� (�$8k�w�`G�L_u}�UWлk�;�����%]�76������)���
# l�I��pN���C��>O�9���1�&������a�H��0�_��EQ�>6���-�24��dv�,C�������*
�Z��.�
���@�F�#�	�Om�q���Tʨ0T��:�n�L�F)s{	�ю��"P=�h������T$��������QGx�����`����"���z�FXd��y��:y�3¦۞���@L�!)+��2��}�����G�����g��V��J�������0�D)����t3b�1�c;H�m�ye�"�A2�B�J�us������a��ii���VQ�	��jT�+1TM�0l1/���v�1����s�[*W��sX���,3[�3E���hwb��,	�T��3��D�0KC ���[�	��bv6~|L�o��nyS@�/�e�/Y����SL�^Iv;�W�6u�zZ:l4B�^>�(`���	����dUm�m�Z߾]��x��d�'&�/z$fCMŔ[�]Q8x���v�))�w�&T���Ǻ^�??��i�>��b�
hQ�=I�g����xz���#{���A�゘^X�s�������v�����<�� ��`�='s���"�<l�	ƛqa�٘�*��Q�]��)���z��0r\�T@�!������K���И����XC�(��k�*G��I��+�D�˅�5�C�=I��ݻ��*Xإ5m�H����8_���c�uI!0� ��P�䩲S"���Ie���E�.;�R�X�ޟG�qf�͇�hZ��#�������L5[ǧ��U��ϯ������Q.�6'=�j�I�_���)'/AC�g����ő��ŵþb��=��n�տA<͠�[Z	�<�]���L>Ѐ��Y+��T����9n~�fL��[�� <�"O�K����(kTWW�H��j���l~'ʺ[�/4 J���/��]m����wo�lu�	ݭdg:;d���^�?)8%m ���.�Ne:���R�Y2���^�P�-@��=&�ƹI>oW`��Z]���0�7a׈��)��\�ո����⟺����G�װ][9��e�<o�H������,�.%����p(���������#` �`I��&Ⱦ���>�q�\��ND.�˫�X*U�.+��d9��Ϟ���;r ?g�t�/]�%��-`/(�#�WU� z����d8NI�
?	�S?�Ж��A�ݲ�X$��X �x������,h�s�a��W;����ԕ��8$��H%����ϰ���R��^t�9I腜�Wｉ���]o��5b��%ݢF�mQn8H�yβDz5��骎B�7����?�t}��Jι��9 .~콗$-� ����r�A-�)&t� �H��A�Uq�n��J ohڷG,���i������� DLBٽy}�8rp�[��'{,8�d"���Ƭ���T�s�k��/)H��c�$x��\)��$�7�I������k�*����u��~g�d�<���G�g]��5©i��xǢNb�B���,�E�`F��d�!oyˉ�}W��/A�\��ř�0_|�3�����m�O��L$� �a�n;��9�F�>�9���~avD,�a������uV˦B�Pp��d��+�1�w�]����r		�tq��с��v�Q����͊�X$$�w��S�3
�����So��W;%�����2Pg,Iln���| ���K�����h�(M.$��[Zh���+���K`qc�`En0:�~��_q�_ɣ&�_�o�.�I�Nڨ%�O�
J|�_h_�/*�j�����~/��E�2G�r�3�-_����J�t��HMXB���n�D ���F[׬B���Dɋ�5*���PZ����o|)�l��Z�t
M�)��i��K��	ĕ��H嫃M
=:x�>4�kb���T�(9�M��k��}H���$d׍_AMl��l6�j��WlI~<Y����M<�&�����KV��6W�
h�1�Ě��k��.�+��H� Dpɬ���$�.8�[W9(�a1�M2،��V��Ԑsg���J^�������jҒ�ƀ�2�4q��^����cJ�(��ʳ�9	FK�������N�8[���e�@=e70����˾YK�rJvg$��b��)�ZE�z�%�BƓC��C=s�`�&�n޺켑��a��&�jnVNQ�5�v|*߆��Ed�W��!NuV$פ����ωM��+��v{8!Ɵ�o��um.��� D��/9�y��g�l�aZu���-x1�/��9	V��S�2��x��1J׬YHH[�x-�µޑw&r}�X#��E�ڕ���.%�`f����f��+8�!��ս	Y�!�>͟���&8�N,�>�z)!f^��P[�:\A�����L̃;��.���:���p�����j�x�pr��Տ�#J�@��ѵZ.�۩����L7�1.����Es�}��=YΓ�B�(��;R��$��,E�)�.7��k��T�y0��a��;�h��AS�y�uz9�q�Xzo�d��slh���\:�ۋ
�bl�5^��Oq��ˈǼ�%��#"��Qz�$��[zG��@�7�%Qj�
X�xufX^�j����l�[jr�$hh���/���L^�֭�`3����������yѱ�%Yq���&��7���$U���8����sw[��-x�7��o�=#fol\�Q��DG�N`R0ǹ#�#ᠧ`����=^ؚ�o	Lh=Ґ�[x&�ϋE��^dl�c���ބY���|�#U�(+#a����)\	�1�F��1еa	O�������PG��Lf�Ϣ������-*�/�řh��q�c5�Ұ ��|l�a���H��r���>?�v���#nlRzN�tT�^�`@��c^�a'���ޫ�w�2g�z�m����%�e�'���ސl�����y��3�4Z"���,��_�v�z�#G����r�מn,L,����R�E�ؽ�iԎ��k�÷*Fw�C�_Ö~F�.��T�dH~�ey�1)�~��Ä��1p�N�aW�K�b�8^�9�q�nb}�R��;�vR�2��/K�ڜ��q��:���8�%����,���<�?����W�.B��BP���4�ђw����&��s#�IW9תŌ2�C�rSt�8���v��J���_�#�rvf��U�8�L���D��7��̭v\iz�8QAM���	<kì5{>��8z���e���:�q���(�LȚ��J��W5YI��KqC��skb]Ƭ���n�"�5Yx�Y-b�����(_\�R�rY~�SN/oT��Tx�Qph�Cߚ�^(�YJӪ�� Щ\6Z��P�-{�f����4+H��;#���>��-�4h�G�̤�~�1se��H�f\ �D����s^hn!��F��o��e3Y�bMw)��j*M�`����Hs�Y�@p�kk|��d{�H��N��]���;����/���&V�����ó��KP~s����[_�Z舴,y�2��k =XF'���/D��F�O/�ǌ�����.�GE1���9YqF��^����fJ��%�]���>��n�r\���rty5)+I%��s'e�a#����UË�V�;�SIG���SKn��eD���)��y�3�.؝!�1��?��,�,`��A`6����PfaD�=1o�i��I�	�۽H�ybF9fX�-4������.pu�Z���5�=�X�ˌ���,��,�c��9Uԡ��>1pZsY���o�0�W�	�	4��*1�����#]M��z�9���F��ʇF�Q���խF���P}�r�Z  p��\��MN�)&{��+��$��Ny[h�����ų���_Ovߢ��nZ  �2����w~`t�!X�`X���������fH�������W?��`B�W*����q]�����߅��N���鷯�D`f��G�2x�6y� :�����k�q(���wVr7���/����ٝ�_l��
1���P�`��?�A$���d&a늳�zg���?�!wJ/�u��U|L:[
��KA�&�F�Y&���;�'����|w'�T��/RY�n���@eB��է�ו^�/(�Q�Ҹ�7J>��6� ႋ~����dw
:j��*�)��#�s0^Z�Q7fhz�5�PG��.4?Z�0&���2���8���/����z&� ��8�8�5B�-�G@���j\/O[[u�L	��8:�2�3�Fl3ƺ�N����ٲ�Y�Ob�O&QTH�Ut��h�R)�J�>�"�.�0���He�k����+�2<�/o���a돿����Pش(����ۡ߃k�C;'I��+a*�JfvB�W�À�b{E]�/_���a����c(������Uj~[]h"�/���,#��eT�췾�j����,�
?��(��fX/��;E'�;!�j�9|�v$Y#oQ�L}0��F?!u�/�Xg��א�A5T�Y-e�_[��qMݍ\ز|���c����^��j?�sg�E3a�w�K]d�y��E��0��bY��ңׄC?���çH��"12�QD��s��O�����~ʌ2��:�y�֕h��*�\6����S�M�~�z���1�ƲE	���N?��4řVK���y&�Pk����y�����s�������\h�Eԑ�D�>�H0�����I4�Ϯ��y��n��#�aXs1�~��c�{E�9B�d����Z>Z��1ٳ
�x� ���l�3@U�4�R%����K��An����]l)o����f��W�X\,泴��h�a���B��j�)&%LVXg�R�殰�� g�dGW�{�d���D�m��?T,��>Gp��0ţPKtJ`�d 4:#KK�b22
Z�z^O�x�"^c7�f����?ɭ�^.��>=�Ho�u
�n\DG���3&m�E'N��
�L�_�������|Yx0	�U�u�q��.>>��O�aUgU�:��X����Ŕ	��w��m�L��vg3⭎S��rЍ����!��nE��l=�#���)E�-�\o\L��Ё'��,�S��a��k�	ԕ�rÏݮ �s�ǲ���+Ic�@E�X-��������K���0�̭��l���{���i�/��o���3����x�3� l����ޙ�^,}�笍�]Qa��C�.t�<�ZH�
��{��efL�?Ȯ�^ܯ1�>ݘ욉-��A������K����:��h���>Eo��0R��S~>K���3$�1�Ѻ��m@[��D���K�e��L��賣Z�m��0��S�9��
��X���չCN�+�-�Q%����� ��d{1V	��T5# q4av~� с���>�PG�S勞6R��/�&p�_�}�e�Dw��x
p�"���j��1u�(�Lĸ�\�� �+MR�-B����n��	s6�i�2VHUw[�ܡ�v�}�W �:�m�����7�l�g�vLP_{�e�w�D��C�WHFQS����Vx�o{+o��C��1s�+0�n2;Ԋ��MP�R9��* 4�S$z�t�Ʉ4Y`�n~k1LR���N>��մ6=(���y��;�nXũ���X$�����؛�aF�p�@���� �|᜹3E�rF=������2O�X������J cc������)�����ol
d�=�y�t�U���e)�\}�s�;G��W�GA`�]֏[�s�����ʯr,>(E�Y��J�3���b���BK��
~ZZ���H��3�9	V����p_�^F~�'�&2���*>����ZE�!P
>����Jg"7o0��D��r���f�t���{g�j4�1-T�ha=�.���4���c��vgr�6��Ϭ���g����ks}������ 	�֌C���އD��ZPMMb�Ρ�e��&��9	��#�8�مf���0��Q|�QP�R "܆� Iv �JC`�}cI��/O��|�x�����Ñ�ʚX���_Y$z�q�� v�i�^��E��{�-��?\�"pV-��=Y�J,���tNl`P��]�G!��*�U��bk�G��Q^���6xʁ�|�����jZ)�ؽ�@O�b����,����Z*J�=���4��v�7[Ԏ7^_���_���yUT:jH��TxT�S��w�/GzG�;[m����*�U�(t�_�h�F���.�|��%��G����(Hv�"$#��Ep��F�S���9�L�fFGLNݪ���.{�m5ej���/=�ʭu`��~���ّ����3��M=|�H�U'�pti"-v#73�{BTM �NG|{����d�x�Tڸ8���G3{%�6�����Lvǯ��BH��O��uP�/}Ű��5O*9!��N.����&=��b�`�t���Jt=1�e�H����/y7sL�5+l���{�կ�*ˊ�]���5���Z��*�����4�)Gz}�[�)�$��y�P��k�G��U��o~
�YYYaQ����k�?�Pk����m-�~K{��쎪��;}���C叕���S�k;WqD�?�^ILܷ=h����9��D���gȚ�EK���lK�>��l�/�𽊳|��Wx���>k ������\��uņA�y�A��-�1r+45%e�U%�� +���.�떑�j �W	�%���Ƅ���c�|W�©��~�^�
���Π���]�]0�y�QCx�"Z9�wEن%�R����qi�V��|�ִ��ՌN���u5�$:+�$���gW�܈�na���G⓮[��q�.�T���ħ����h-\� O��M��&�v Zj�z�x��3���ODJ[rb�f}���;����I�/��f�����';���.�cWu����h�[R�_{0)����9�2�P]�AZ�O(���G�Oy }��8��Vp9���	ƪ�U|P��;CW�=����be[��oZlah\I�~j��MKJ:��D6��{�ߴ��}��H@09�C���p>��9��T���v~�
6���r�p܇)��9�~��ûp#�,��#5d~�������c
(��o�r5?7�>�F�q�\"jlL���C3�LxL$�AGkC�Nl�^%exc��Sș���I} �Z��c�RY5��4����i�/���sͱ�wAY�V�fK��l��hh��J���\Ȕ�� v����/����G�Cs7�?�+���+eSʬ�)G�U�u�4"��ZO�@�(5�_~�9��e��]	
�����d�	ubA
�=��B�^PƓA�������4p�
;�:��"#�~���L<��f��7�����'��1�d:b�̴4�)���1W�����P9K���6)#����1����hQ�E�7��=�4������S��][����h�=��C;�����3���k��z�4��`�s������&s	�q�'[vF�h��,V�a�~!K�/���_�F�UG�������O���, Sy{ �5�̸�jZ�ֻ�[�5���ܑ�׋��3� ����b^���73�R�#��0�Α�����ڳ�e��=���Cu>u骭ɮ���#i�ñ��ǳo������ϓ�\!#�����U^!(�%7e�\��mVi~lؗ����(@�U��,�x9N��UF�'S
��"��۶�W_P_�\p�ho�' �v���
Ok�.ύ�
 tP���D�"�w�q_2�fퟙ)�]w���i64=��?��Q�RLX���r*�#�F8臄cT[�'i
������UDϩ�S+��a0l�����Ӂ�ʧA8�(�RҶ�y6SA:d�d~WăƼ�NV4�T�ҝϷ����r��X�*�^����C��l|����K���8�(J��a=�mՈ^�@����#�����L�;T����,����oݤa᳗�c�2���!�K�"�����^"A�����cK�4��;��Q��_�X:il������1yaeEV���zx7�+���?��v��Bf|#N��=��H(�d��ZD�������uP&�N������_H��軒u��8��������,�y%� t�<����vM�_���͔�ݱ�����I�&�+��vI���\���I-hAZ �<b;��CC�T��*���@��u�z�u�O�{w
�΀�4��XͿ*\��iVlRUBl�&��4>N���ϥ�����\��@vK�$���f��x�,�p4H�B�c��k�7s:��v�H	���82I�q&�W�^�6�9q�8�E�^� ��L�b�)|fQ���|�#A&��C~�9�U�Ɉ�W�I�����2��l	9��?�Y໰�N
�����s���S�s���F*I#��7���/�9�U�k�-�YgO=�ҩ��Q�Z_*C�ŏz~���D]z���hj�S=�n��3����eA�$�D�T��i6po(Fqc��PRo>����KM��@gXÅۯ�C�1����-��),�#�1(���ƃͽ-g�)0�Lʼ�?���g�f%ʷ�KC�(�[�Nw�a��
�;_�NGB�T�<H=7Ko�� +�tw=�֪�/�+�,]l��*���.B0j��.��������/�H����$��NY�|�w�67� +_y������=_C$,ܜ���!���]i�o���~ks
�=�-:��;�D�P�Ai�yM��YQmY��#����TEe$����@)��O��¬��j��s�j��5�H��CK+�[��%���D���Z�H*7�������~��w��S���٫w|�	X�yP�O2-�"�B���Âj�U]�������|�C�ԟ8ՆH�D�FT�`�YT7�Z ����� �]��2�#�[���o�ǈ"z�s����tn��\�z������irw��8���ժs�jJ��`�H�j&���R�ɹ>� N;E�3{z�#5P,�q��B۞�䂺���x4A�g��W���5���g4p�e�w��`�[JC��L��ٳ'�\ou���s�n _w�g�7>� �k<�>�5��81�i�K����ut���C�w{��Pf�q�o#q#�ql�l{5���3�=�Sw�"�jB#q60⣫P�L���'����2�t��w5�V����=��+��Yd�&Q��x՛�S�dz���>���|E�7'.��z9�	e���$�: W�L^Ûa��>:}���-�5$��E'�?խ�wW
lJ)�k�}�\x�p<A7K)�@��f̀��$�(Yy���* 2������r�Vメ�/�p��S+#���};�&��s?%5�%�Ěl�'�p�,`�eL�C��o���_j]1��k�3\����.�7Ì�\W������R��`�~P�4�(��h���j�
bڪR6�3Q�x�����D����
g�#5��N�ƍ�lp�����r.~�����8 f�bԳ�*��x��m$�J�=���Y'�#f�y�� 6gk�y9Y��o�Y=fĨ}ֶ��J�B	$�w�R9S�(���g��|����� �E)e+�������)�����]�D(eN4AԮн�P��x�}!��iV�;,?���:��}M��ו`eROq���>����5~�p��!���m���N_r!P��K�)�6Ϻ�LP����4'����rh�G��:����W��Y�,�Qe�#[#����tpz�dI�� ?��A�9^s�o:A- u��ڎ�I�X�̩qn����\I4���~꫊�]s�}��X;�́L�?&�H��ظ��_����TO��J��+S�EF"�7��5�V����롌�Ӄ6àӆ�v�˘j�S�8��S���1��^[3�DT���/���
G�X�1�_�~$@s�2�����?8B�a�N�S[�����CA����FQa��%��5�$c�V��z����ߴSnޏ��1غ�9�0��o����i�"_�=��L|3��7�ڌ��!�8B�g���Od�sd��|1��M��ꐞ�kT>`km.��u?�����o�bS�9E���~U�j�RG?@eѡ����im�.��;5��, ���/�*�PO���`Ɣ���ܖ�7{�G%�����C&�8;:����e��̏����fO�lJ�?q�()
�7��c
өA�T��;zM�'Rq� y=Ѥn�}�e�6H<��@�����м\
JX�|��@�6����B}��
�=�Q��,67 e[U�k��������&a`�#���4/�E6\@��3�x$}�sd���&G�c��(d���$�զ)�껿g���M�F���j���E�r!n��f���d�+Pdj��`v��C%�\���ŋKկr�c��Y�:����e�$�l�Ǵ[��s�o ;�e-2��B;��Ɯ>LIwK���"8���	����%ԛ����ӻ�bV�E��5Χ/E ?[�UrO3�1׿��xob]pGp�}������>s� �A8n˭c��>���AÐ���xֺ�s�������G ��r�CQ��V���vd�5p��"I�[
��n��X��

�<��wU�[�y�/Fڞ@(�4V�#5��q{=CED^)���k�CE��^��#��?;ݔ����j�v�H�O&i�gM~��⧯��"8����ÞY}e)5��d��g+��vqdc邪S�"��r�գ��U2�t�n�\M6'\w:*�۪�"a��+l�Rj�<�5��2��Kw�R]`��9E�F�]��⽄�	���N�M����Z'ĸP������3�߀���|=6��5�v�o><ҋ�Lx[�J��Sҟ�*3�������׍V��r���LY��g�-������RlCs..\�D�ʊ@���zuϝ@"po�-p�\���G�7�1�m2 O#�YM�!KR֥1��z�{?����(@:��_̒�1)�k�*����>l���f�����p�L���w;*�O���;r��O��J���]T�^��>9>�I�gd��j7N�~i�:��첖H�ZH`�
�L#{{�Y[�OsL��D=熎�'f����zU��w��SfCju����¡~t@5٠A_�ʜ��J���<?K1(xIv�?>�c�#|�\h�(~K����+���N����S�����C4�٦ۢr��x��r���1T���:�G��
�������
��t%\G���M���+��Z�o_H��i���=@`��P�o��n0���g���{���.�_�f�Ƅb����z��X`t�s#w�s^M��`Gg�W/t��y� ��20UzV�b-����Eq�5̌At ��k1!tV���p���%����#��r�N�������#�;q�3�J�_�ݡ������!���� �˫�TO}q��9�,v��3�9@���j��4�o�%Up'"�0�[B&g"Z5 �<=,�1ˢp� ]R�i,�=pb��P�1���V	B�6����֝ҳU8�d���}�C���1A��7\�Ԏ�c�o����x&���#W���KRW<u���-�`ګ��ؒ]1��Km� ^ �k���9l�	�5'ֿ�3��#rO5��yݼ=�Ms��0�I��r��h�������.g�a4�m�$Dz2(�F%��\���ҋFqI�m��H�EI��3��׌���'Hl\Yv5�^�+.�D����d[����|,.]�V��yc�g92M�2�g��JOׄ!�������Kg��H�>�Qt�Z�7��q�k�W,a_�G�5��QmZ6��roF�	�V�o�9�넹�E�O���	v�V���ޯ;PbS����(	�܇�S{��d�;��#c��'�ck=�|� &�J5ʇ��Hu�3��h+�55Ȇ9ƹ@��x�{�nx^hVi���ؘ���dx=�[��?�d��+-d���.�+â3�^<"2i�M4
b����-�l&���e�2b�G�mp��Z8��N0*�Sx׬h[-ɲ��*��k\�N�K�cB\����;��&Dm�h���yP����_	��F�����n��TwϢ�&L��j�jm���Qz�4PL���Z	�n�vC3QoX��9�����p���D|�Z�%A���TF�St-���K*j̤&� �]���&=����g|ل,����a}VNȏ����p�:�)�T��꽣ՖQ�wAM�Q���V�|�92֗x.<�T����?�4J�R����h�٤�H�_��^��[P�e��.z%�詩���f�|,�~p"ۭ]���Ca����	�6�I��ӣ�?ՕG�v��@�#(�ڂ�	�c�����'|0��.T)T��Ϊ�Q��y��s�G�b�W�e���c��P�[�=P`2H�(�Nj��K�V���-樳���b��H�=j&p���a��9����ز��H�@��Y9/�UjJ͚��9qm�8�I���j��ʹU���v�J��YY;��п��\�P��PRFDZ�FR�n��E,��O��p���"-����A_>�9�!���`�!#�����=��2B�%�3���X-Z��H�Nډf�cQw��[��B;t'mɋ7�\���ȼ�
��hs���	�^R��N��`z��i��GhR��[m� �a�R�+ӥ���H9���lH����xA��P�^�����$L9=7�^*�6"_"J;BS�F��6_8b��'���X���ℿ+�q]�~��3嬦xC�.������ �����\�z�U�Ai����	�I�[���j�rD^�	*NLC�B���nN��.sl��P�qȸ��_����&����e�r9���TW�bx�=8����3�	�(�m+a���:�p �:��fq���AIi��J����#&�b��6ة��qQ��d�8v������{�B�B0K�c�P9�'�F��m$�����\նq�1F�F���&h3
ڻ?�Acx��c�^��T���&%Xq-��ޟ�T����'��#�;�����(���g
����ԏR��'W�,����"����mrAäRdN����]<�N~���8�\B�1j���y���,"]v|(�&!vA�3s�5�荵.�-�K�c��NXk.����W�梀���q`n�^��cAm�M M{k	���N��8���)��F�T��i��1�[��������+;F�@9�9�Æ�0p�ُ���
W��ˀ�M�{<��p5U��ơZ����I#��e4~7atg���ӑ�h���*I
d�Խ�qq]���H�ҩO������0���hl��ʃy�@��E�@� �C��[O��yJ���kP�S�W��=�5;7(81�k�4В���U����ܝttqYΪT|�(������|Rh�q^�M�R��%]��A�|���X�;@t�F�!n��;���\v�W:h��66?��Om���'�XG�2� �zZG���w�2)��C~���k�R�s�b u��ēZ`�9�/7�a¾"^��0�x��)��{<���-�ċ��ۣ� +j<=���|��Bg���7�*>���R�H��l[GdE��� eJ�`�VX�2?��%������E) åֵ!���� ��TBk�o�mo?ʧ�]ۅP��q���V$���A�'��7P�	�o������AcX����jD���\3Ʊ�����&3��j�e C*y��B�p>����`e�@1v忈R&P#&p�r��ǅYE�ּ�{_��9������֍2��J]J	/�-��Z[����
D�(e©�������e;gqfb�n��fώӰAٗN��u\�~�)5I���'��g�`��������	bQ~/u%W)+ߥ��h=���=x�Rx�N��c�o�Ym�	�}�w5e8h�tkZ�@�����:nҊ�Հkpu�dW��56��.��K�tw?����t���u�c��Z&�W[0!��Zu���]_8^�n�X�g�|����4mn�ڪW�.#����ݽZ�V���-:M��f��?��B���.�wv�_�w5h��-�6�uBgˁ��F�( 5�0�b���{��{(f���O�~���iP��_���U�����[*aޒ~�(#�_���xŒ���L�uҽh��cs�F ��dR�)��l�%�W�$!{:gHBf�}��7�bN~%����[Yl[t�p��.�w3�5����P�B�� ��E�T��g�y�\8\_S�I2%��/= ��Cf���"�h�_�,���,|��2�{? �#�����y�I�MZGp�PȻ��}z�/�u��.f嶿k0ZQB�.�KI��<�GG�$6z��c�Ĩ5Dk��1��Zh4�{��|�9��6�a3;���O��S�J��\��[�e��@u�T4�8WF��UXP��Mۦ��^m+���i�5#R���5�#/4V�iYE/`���B��JvLz�&��|��>P�5�4 ��f�'L��%>�U;	�������m-Qf���
Y����!M5���Ѽ4��qj��*��`���)���l{�+5�6�Rym��E��|�#p�r������L�2�{�+Gl�Xj�����]>�Ю=���QCi�C��P�6��%��3,�����R~G2"@Z+�͹��-���3Q�q�[n�F��e��V����n$Y=��z��ڸ��f���2� ��^�9����4V���L�$|>
jK\�4$��3ԉH�(��%\���a�/��nk����%)x�A�}��@J�T���Q�����`�U�6�5+ZU��Ȏ��08ي[�'X���X��*F����L�=�7�����ch�[F�~Z�ZÇE"��ң�#�C֬/��S�؍�곛N�ߵ�7�(�F]A��Wޏt������{%�K��1}����Z���|� io��l�VI{L�ʽ�X�?�3Ρ(��tw��x�:7q��.��\g�a	� '�3�'�-X��T�|�I���O+�e��1B갖���e�܂��\Q� a�����g�B���8F�j���Lzqm��֊��e'*�t���*-ϝ�J��v���0m�X	�2E���2>w�3��'��w����Fb0� �0��F��d�A��4��WOj�d���)��UU�H��E
<}��m9cS?}j�F֤�OM�:������)(��#r1�����u]� c|B����	�eS%��H�ѽ�.���"��5
ϴM_lVƹ�~��)L(���� �u7j�p�3B��/��Ӯ�)�;�W��W�3�e\��&�v�}bpf-(A\SIg�
k
W�t���:�O�8W��˜��f+��%j0�'�#�:g'�{e�nE+�k���A,$;�k�s���.;b�ޫx��&7Ts��F:����%�W���*��ĈA8�Q���4Ǻ�0�aQ��^�,����.lmJ��0�g�%U�ذs���s�&��Yb�'���&�������%)�p���y��f�p��B0�W���a'{��A!�#�������3o�y�zX�K����N7]��T��^S[�4�X�0�]�:���Lo���z_��y]�P�>�`
0����dt�6�5�0
��b$$3?K�&��/Ԍ�������<�xČy��[HO\չ���������C9'Ȱ-��ԻK�t6���k6����\���_����ldݙ`��M~p�,��r�;z&�-�'�s A���CtJ!_���2ݗ�W�a%#����s��`����������.��u!>��_'�7�mN[I�)����O؊��ޑ�Y��A
R�W����x���n��5_�a&1�{�(8٣��<�9vXz�z}w�7Q�Pl��1���~��h��yH�6w���a�5�?��98X�mHׁ�s���c�����?��`\��=eIz����8�kL╺h��f�;i�kE?�t����u�ʘ�?v�j��eo������#&��!���R%�[�|�өU"�e��YN O0��Q���*�(ۖ���Kd���2fsG�aXʺg��b ��T�8�_DRQ#GEEY�w�[*X�8�4��(h��J
����z.i~�:�������^���
��P~��C�O�H�Q�#� �M-�Gi)�-.#ܷm�芿@B%��W�ON/�������F?�?{9"�d�A="���Sݚ��]v�\'H<�68ss��@�d*��/յ}~-���������nl���pي���0�o�S���}-���3�b����af�2��ň@����K�Vä�2��\Ktv�mRq�ƐmyR������S��W�#�׍�M��j?fS�Dph&����sv�6%^��G��T~)vb@�2��x��RV����,�&u�����gD�)����
.���9�!~S���:W����b��|�d b��	ӛ����B>��}L��M�%>���<����d�����d[�,-����>6^��+P�"R�y��-&�6V��e�.�T�X'���~'����-\�&�j��Y�X��h�DD?W!�	��.�ӓ���iL��������lߦiUX��:�tq���n�r�֌{s����L�K�� ��|��FY
�i��X�Ec��If��ԘM�mm�vDZ65��VTe���$�&�m�jq(���Ĳ���8���H�t+F��c���<܇I���^���ԆDB�t2a_��$��N7]T���Eê~��$֓V�$5�t�j��h�bK�8,\�.�kHFk��mlFD�m����2�l7�J�U��E�2®8<kR-9!����j�����.��x����{4��3|g�����c�碌Qy�ٺRΆ&hK-��������GmPf�{W�S�|X�\�\w=�f1�
�K���Y�ʄ�`p�qZ�u������	o�1:S��Ž�i��i�s��K�uZ����KH�������	�M$���e�	y(2<7����*+��CD:�k���Hͨ/����"(������)�v
�#o8Wh�V��$wc���_y�sq���g��:YO�M� ��seh��0mƨ/I���K#�x�D�h&i�oEӊd8�"A�2��� �D�Rq��&�Vwۨ�Fa��f�G2E�BL$�RL���;���y7d�*/߈,����n��@I4�mX.�9���O��O�5��<�dl�u��`�Q  ����, M��.��09��^c�Pvo��X��?�:�t�}��⃁�A�W��ti����K��}�P�}�XQ������&�/Q`��b�����EC��v+5#^��U�*�a`�� w2�vI�_�EL�$�u�7��óGp'SiӖ���"Sm�"�K�_���E������� ��\r�?�����Z�D��*��!5B�Y��\R��m*@��[� �@��)��iMñmL2s;�<���$W�O,�A�Z�c�܄V�!��)��*�5G4hf�W��	�(��s}����'���H�r���w��4��r��Ր�� ���u7�LC�8��nxHJ��NN��Y�>MRa�Ǒsep����#í���D��yT�Og^��P�{�X	�m����f�}D�Z���f��&��c�A��ϣ�\<R'�i�g~��Q�K�i�8��QGr@����,W�6�ٛQ����'���*�c1m�a�r�XA��D�3�<d-&PW��$�mPF�z�n�s�l~�N�4ʐfªYt����NfS�C�(��� �)OO���b�$�eZ4�����0V(Q�xx�>���d���U�����6�@U+}y�	C�`|����9Ѿ���=�$�U.��(�꫌u�O'���߹�Q��ߺZ�X��O%h4� ���m�؀�z�NaUp2�}�:A<��߾FS=��DI�m�:l�$p�@�4�J)=�`�jwo�<�/:�v{���nl>�&��o�����Vk����2�T�����<K�	�'I�$4����6�ɢ
�p)�4.>a2���p����AY����;GT/��,ir���!�`�0�kP����Q�|�V�@^��r����6�'�xNN��ɚ:I��p�����1=�9�/bǰ��Q�;4���x瓥V��<r���K��*����G���Q�a�>`�Ԧ�ZH��5�p�E�E���,�!���T�{&�CB��TEV.���4��푦�Ġ����s�/�Q����	���ژX*R�'940q��DQ�Dx<���|f{FJRx�Z�~��n��1�3�����4zj;�������B<�3�P+�dYU\����8w9��
C��S�e�9�,��t��~����R+��SJ�T��ѫJ������菌�p<�FWǸ��w�@uGl~x��j�j���x����<A�.;��r�����/��}9E��2f�l���U�E�TZ�˂/8���k6��Z�(u�i�u^4�Y�B\�>"@���@�~MQ��t�o26�@���-�;�BT����Mb�LM�N�~���? 5���A<��flh�u�	Զ!�wy�?_���H�1sPq�?����y��drG��f$(5|W��|��c���[6�AQ�ʷ�ǉ��NW�Ǎs��L�6;�����Z7jM��M�qߑ0�G�&�ݖ�T����E�u�U�'�!�𦊄��ϱc}M���&���tb��>�*K��#��R?Së���t$��h��ܷ�D�F[,�G:������]�[Ӄ�DS�|�B7��F�-7��eB�H�~]�؝�>�w'c�wH��4��U�J�\��d�oƕ9w�����N1j��bB����f�6��:��G0Ȇ�%r]��n9H�e�r�>���۬N�Qz��[���en�U���Pw؜�K3����'��T��$y�	c��d?��MC�KE�ܳ�*q�ބ"�W�Ɠ���.�@�+�׋�� �t�����ĄCPC cQ���R� f�	j�R-�U��}��>����h���7M�5�ޗ�>�ۍ�����!��:��S���/zhz�ϵ�"�~�ՌFPY�~�;��=$=�x87?T-���Cz�x?"����A28h���%-����'��Z��W���V|[M�u�q����OV�/	�x���6��r`
�1�sD��$x���IͰ b֤7�[9�-{v7�9��1ֽ3�Ê8�������t�Pt��'Q�:aLޤ����&����ĳ�kʰ��ֱ�'lJ ����խ�"V��X�WOQ~�\Z�jΕBW�ݍ�O�\]d=����(�쥼*Z���R�d�{b��=��h�.f]����;9���K��x�Lr5�"wDӋ��0�W=�Wԋ|���}��9���=a�!�,��*X�4E�?l�|q¼}'���~�Uhy����rݼc�v��'���y�\�M!a�37�޷+>�_$��=ЯǃO�9�H�dX_��xxC�}&���^{��C���K�xq��fl��\��A�L�)5e�S��Єijk6Gi�c��GC���|���p�,;���wjV/��(�#{���W(Q�:'��"��j�/a����s��p{L�j�B�����܃�B� ����vD�x�]�Ҧ��c
L���D���$8'9cVl�>��Z�g�Ƙ�`��r 8�.CX%YHc�@�L�2�`����.�棭, �0hʍJ�n��=����a8���kBp�
��ٽ�x���J;h�K�U�Q&0�8,\����΢�d߬���C�v���
8R�{sZ�=���(���?�S��U|�#ٓ�K).�GH� ��T{��aێF��t�H�`�mZ��U��3��=�S�q�(c��|b�Ig7mjF(�� �K��~�M�շ�g#���S����9�j���axL"(�6G|}8��:��9�ΟJ��j2��9��z@6�/Ck�&��#q�>���`	x�zU	��V��<E����8�}�tֻ9���� y���L�OS9p��e���T�/4�A��p��'QR���h�"kE9��y���:Hd(�y�7��Y1?Y1�&�Vf��|�/�l���*�����jc�U����p�(rGCM��v��
s;��୭;? ��K�ޤ���	�F��0�_�-4�uk<��߽�� �8���
9��R�y��O�n�>y�5Y��%���u~��/=6���r����m:%�� #��67V��N��av�-�uF��Z~f/@��E���xetĊ����FHVB����uN뵤]J�f-�:����0��DM;^�9�Z'#����Y���n8قCn]%Mp��ရ���R�6v�����oLAm�>U�TPs/��1RB�J"�i܍?Ң����lnCh+x%���7dS=���_��q~�vf�D%��L����[@-k~����8ڐ99k�Wl��[�l�K2���M���v��]�$���{M;�h��:�`&nsTk窂�{�81qa'�8ƽ6�&�'����d�ͽZM=!M�����S��"�����W?�e����(xӠ�� +��>��F���W��S��T��Ѻ���t�<
��vwk,�Su�����7�pz��{�lc:�%@<��J�z�dPP}�Z����c���ղO
��ռm�kB!4�<P@�����;�E��ñ�K��.�N3���]�Г�6D��$�rQ� I�CR#ˏ���ci�=���2}�f�>���[
��`��e��w�ƍ#��gg�'�}`β`�n�|wIS��ʡ���7(�$����@�"3�A�r�{ �x���-GO�h�	��:��ʯ4�k޺a|�7��K?7��dj���j�85�_96 qÐv�ÔҐ`���9sv-��ۑ�!���P�h���O����y�Ԏ�1Y��n��Z ��6�Zp"�����s�m�X6�Y���4Z�&z�w����ݐ�(�x�8V��qT���q��-��Q��2�1u9�}{�{���ԟ�H�E�S���ʝ׭<�b]Bg�S/�|�� w�-�:����!g�|��C�kuf�U�̯-��O�U#�;uc�wV,Îי��-�/�e�R�l�0�~W��5���y��Q��6���I��	�����;���/(h�G���è\�qby��ǉ�RK����8H�_u�*D��(O�.��%�����A�qJ�F4�	m��ײM�2O�nIYC���4�A��a��B����7��2�p�G8;
����(��<�P����k�{,~�x�5� �H�lW;���7�,��}<
���pZ������;���&���³������D����6��YǬ�>q�|�o��2����%�xLt*�M�� Q�[��Пe�4{]fwH���@�%����F雦,�{N��Ïo��#9�4��#EsA&���t���`�6*�ū�k��S[�U{�W{E����Zq����v��Z��}0y�( �\��$���o9�W5RR� �U���q��F���,
HQ��a�c�CeM�R1v���R���]��F��;�Έk�m��#���
�Y�k�㺐�2�e2����%�&f�2��9�E�qń���Hg΋��m�e�,�K[.���`��yH��U"��فo)�&��S��0p�uHY�C�|����hї��ᭇ��<G%���Ӄ�pS��D��)ꃔ��s������4�=�i�yd?8�z�ObQ�}1�~QOԘ��f����o�TγA��W�>,MgC@Ť߬v݁%���C��Ȩ�2B>Xм�J�f8��F$��	�����Aa����d�3�VtD,��E�Kx`�e�w�Lou�I�)��.���S����י9`[���7�����T�{B�pt ��i���;O�����6!���j�s�ʉ@��nT�O�70��)�]��X�#x+���np���T��*p��RYS�?�G(H_�aC9WO(+�o.`�M�*08.�X��qy�'"h��L�V�*+.��$�l��� �6��|c1� ���ѭ�F�8�Qmv;�y������F���Ļg���Z<`�K�"lFV���8�����2��vZ��zPx�apCqĢ�N�#s9���Fe'���(��dX��^��b�1��������l��0�)2��o���!�J��</����V�����x�5���.FD ���;��-X��� �NV�f��n��<j���T��f���>懟Q���O=/^�,�(��1WN����G�������va<��*�X��	��1��]�Pah��c�_����*�&�7�Lms5�� ���Ս7���b�@��!+`U���B�o�y�ʳ��z03�{�`zj;L���(g�	�\�0�RߨM�~�f� �*[3���☉Ip����a'����4%G ��虔�x:������	j)��1���T������ͣ��e�ߜ1!�ߕ��C���N�Å������^:\B��	�1h9W_d)Fuj�[���p���7��(��-X��	j�ӈ�Z�A� 8�Cx݌��M��KG3)>� ��q�pܻ ���>��6Y|1����K,t�ž�
fN�wx�w.�S[5�l�f8�R*Lzl�2N�/�UE�uAME�{85e���zJ�-�t�&��������ߜ|��4���ؙjP;��2�P�qO��A���`����t����K�=�:U�"�����qJ��w���TK�����(T��y���X���2��	:g��Q����4v�|�#��c�𧰊ײ�����jn���'���,��|wί<�2�sJtx���EU;�E�6�)��(�2%2�뜪��sh�`�7F��wx��
�&���o,h����6oNh+����E�`���A��F;ƭe�C�J��|��n3���-Ђ���A�qVH�GD�3���"Y�$`���gR�n*$�-l�?G��H$��3�ng�_�=OH64f������$M#��6��m3������*�j�˅]���QJ�C�62z
�FB#��t��q2%C�1��P-w���Bޔ��mQC��;"�[9�K!��
��e%n��B��fT]GO��Mt C���)H\A�&�J�����������q�g��U���kEc�Az�$���ɠ�]i�����l;���X:Sc��)�̌�5Y�����P�@?���<GV�����c��l`1U;u���]7K��a���1�l��N���b���ִ�	�='`�������P��gL�+{�3s�Y��#��y1�OSH2ʿgn�ȳ��a͖l�y*�dבE&o����PӚS�4[H Z��GR �T���ʎ�yfX> ���\��p�=��������<J>��
���Z��W>�t��J���#�k,t0ڒ��_�d���c��a:��*���q�x�'͚��UD3G�����X��ѱ�CoXpc��&���"M}�'�9��P(>�?��1�_1�b�w���_���|$��d����G3D�l�����yy����"�/rB���=�,�\���1&��P���!G�/y���mźIU�e A� [1uq�1vI�<oGR�]6�壔aQ���,-凵*T�+�����qsk؍����cwe�X�nv�;M�B м���Ue0��5xRd�7
>��������&7)���_%
�>L�0֟���P���;���U^��{7�c�o���h<0#G#3?�o��E
�_t�2@�,��\qi,״;�|^�<�(��ĵ�\\�9:b���x;1[!��i{/���I=�I}C ��s
�-M
��dnqeȲK`�>ߒ4�iᮈ�g�]���\��\�a*����^��%w�C+��*w�H5F,�R�m�n�����C�ղ�͌l����*�rS�/�"��?S�Bb��
>X��=Ȉ��֫C��9040pJ)G�f�l��	��"D0j��W&f�23�?=<�H���5��*�x��;��찳"N{�^��l��#6|.��2Ў�uxMC��,4��}i�c�+m�ľ�Xn�D�b����R�n1/Q#�k�_R)u���4�	����'�(^#��%�KX��*+w�%�@@��y�hAdD�]�C�?<�(f#�����|�rM�c>�����!s�y���h�1�:�`h7��$�g�,��d�����z��_�`�)��D��^c� Iu]~�p|�'})+Ze�aӫ�{������"�b�d"b��!H|١t�䘁�ީIQ�$�(ܠG?�=��%`5xn����忼o(! 55/���'c氼�uU������W�i�p�h9θO~#��9�F�����1V�m>_,��]X�������2�	���Ü�Fw��Ou��M60OQp(Wa��@s����{4fZpQM�0m��O�`�*�����_�у�1��:/ d'2�0v,����m�p8�綔��&�Q��;�%$�.�#��vzDNI��I�I[���Q��{�9c2�O��CI�aSQ�~��Rm��|$�ԓJ��f��]ѽ�yqR���s]9���A��:�]»ֲUd�,�H�J	\ �|��Z"�q�G���g
v��}�!�(�vA�՝G(Z�u�!�ar����#ٝmʹW�d���C�QB�(��A�q��2��p�7��������Os4" �7��*̈́���a�^S��~��4=�E�S�`��RO	xy�b���:� G�(+]`4xb��*s0]!�I�C�tW��U�qYC�!@��@�LxP��H]T1��R��$2]��:��(�3��pR��V�~{�@l>�<Qa<%��~��hܻ��`��4ub}�G��5+gV�pnus\7�E.-���«�r1���$9D�~+#��z�h�qM���O����A�R���S�|���]�E�\�$���5�o:%yUn���7T鰰k���ᛍw"=S/E�)R�S׃#`z��LJ��`��N.B6���f~�ء(}d��V���3Nr�ǋV�6q�$��[5�d��2�Oo����p�d&��}�%�9�������T;ϓ^U	f�Ϻ���$TҤl^}���H6e���~vW}x����Wg�}��~qR^��0q� �[�-��� kk ��_����� ��h������~
��?s`��69�@��F��h�>_6B���,S��ڑ����t���&)gn�Ek-�v�;�1#Ƚ��j�wz�d�^���P|xc1��Z;�B�
����^�[I�
�*z��Ur%0�Y��\��]��g�q-!]���j�̅る?�����{@^�-P���0�`��a\�d��jQ���I��j����R��H�9�%���ӈJ��0���2f"ǲ?	�1�Jj��_sӼ�~��gA�5��(=�S����\#�?�ؿ���I��e�rh'��|U�p��&�2[h4�r����w/p��t�_�\���!`}�|�|��nF�CK�{���sG���M��m=SW�/<�T�	<?��X�W[&V��]��`�)�(��8�Wn/��S�4�ʸ�:@�����4tRDٌ������d~M����Jp����sF����|d�_�:R<��nu9��/}��c�����ސQ�%u���K�j��F��V޹���uc��T���G4-H>k#��}��f{�����㣤�/K���a5bK�!��e^8�Qɝ��z�Co)I��k�?��e�J^��ڨ�U慡�1�pb]IXY��Y˺�Q�ҩztY�L�6��1����d�c2�0�L�H�kИw�¸��Ǖ��V?��VI"������͖��{S�a֜f9o��tt?�X_a��ÎH�89w��=Vob�ߗ�U�O�����>��"����ӵ����ꈙ=�d�Z���=���I2(�|��F�b��*���qho �MQ{��q권�[	�^F+F��L��뗭|#s��d�O�ge��4�h���+�9Ch�������P�<�:�<te�'S��&Xk<�T���~�u��óP��EL�o�ݯK���L�x�^�蔢~Ӷ����{�v;����V���[ �m�$�C�����R�;��];BO���\�1��R��&��Hg�n��殌����2���8ˇ3;Q.�����D��弈:T�?$c�$SQ�����M�����p�@F�h��;�5�g�ז|*��,)�[ׇ?��:I�^��2�e�%���(f%@��"e9��+�HSG����;�|}��^��6Y��܀a��T�we�m`q����C`=�D�Ȱ����J���G�Ƥ�6��4���g]+��^�N� |�A��r�ѾJ��Җ�T��x^9�d�s����]>�x�?tX4go\��� S��0^���7V?�ʀ���Vzㅷ�/"B�3jXEB�,����dWW�s �Ĩ�<����K�j>�8�����H�[$S��@-�L��N�#"��!�1`?0	��x�����iOD�p���FV�e�����u���J�Q�?<D]d�o	�̄�?R��@��^�㗏���d'���Tj>F`�����!��{L��3�&��>���hw3�hk���	�|T�����3u�'�G�^%�0�]�&.��}k@+���ߏ��.��߼�>�5 c[d@���˲�M��a�:-��Ȼ���tJ��6�s- F��I�#k2%�{&Y�L�g ���p�r�}Y&gI�>|� �1���9�g8��40h�����)FZ7��f��p%���D׈b��V���J���)�afK��Jk��W�8>smN��I\/s�^�{5 �f��[;�4N�"z� 1��|��{`»�?p�e�9|5Re�w���|;��2�2���	�PUL���|M���G�S�0&���? �p�/��G��%��ʝ�X����L�BJG������kX��d����^��ǲȁH����>a����35�8lt����c�S�/eP1j�\U��(���\��<s����;�g>�K��hݵ�Nd�N��A��_=1��~��q�7.~}OJ�	�����|z�a�k���qFMyh#=�%�f�!Ja�xJ!���ݑ	�THF�?2}K�M-`��L) �z���~J�;�wJ��-�c�t\8���X�Z��� \��������nr��̱�Qbe�%�,�ٚ�=k�))e��˚Ě'��5)T��U����=/��X����s%�M爂���O��n�[?x��<��2[l�6G�Y��Ej3=�%�Fu��=��L �O�/mY�X$_���Ğ�tEQ1-���?�`����6����](�x7���[l���W>�����r˫P�F莲��*sj�k�px#RB�~�h�*�6�ᠡŋsM�o�ס=d�Ւs9�-Wʙ�p��arȕ�pr^ǔVS\.8c^�t�Z��2*��嵝���[�9�nI����M������N�o\@j� �C5bw^��+��/��¤���'3�J�b3a�����<븞Ä��[��:�W#z�:=Ɵq��+��MI�
Gz��x�����L���P�pc�ΧO��t\s�#o��
��]CI��c��M>F�y�U/ {��4&/����tm��b�� 0�z���T��
���k/j
e�׏�e1��X� j�btU{z#?WM �
A9���~`��4���[��Z�r�l�?t�X�^����h�KfW��ңiC�}�R{XϪA�,��ۅU�{��Ğ�Jpl.�Fs�0�:�BD��7���\�^��ֻ>�8�S$՝׉��dY����F�]��c���,�=U�»��������������ѡ�RX"��!� T%�\���E�%܇����28���n�3���!��,����־���eR�tN��A>'֝/��	�X���J�Ҋ�l,�l��;ɐ�eы�R���RE�^��4�s�vo��5hv����"���Ib�)�|��$b�08�st�k���7�>"���"u�+�i͉�n��Y��e��Ԕ*���!�a�-#'�W������Hm;�%�	��piz�!s�Eh㲙f��X���K�ƻd���MnQ�x�0�)qs�g�v�~:@����*�v�<{	����(Wf��^�f�^�Qq5Gߪ�Q<�֥K�v`���`O<��PHh'�م����{,n�{1�M�x��	���g��R�@7#�����w���'�> �	cj�.�� ��~,�#Q����I���c='�' *79o])������:�F�)�U��XD�!r^��꨻n��|S?��jeSą�Ѓ<������#%���W�u���1(Tl�X95f���,�ޯ�m�h�4:W�H��S7�`Ļċ�K�� Å���e$�}��ŷ�]�JXf��n�x�7�M���ď�D���N����oa�	��9�!��l���o��r�xMU�	�q2#���3w���8I�oٴ`	�P퓝10'�[�Y@c^eŵ��[nl{�d����1��"
U_ǰ���,PKǭ�!:yU��9���yk�=Z�v��I=y�=�r
�/P�6���E��hp��5%��ֹM��$���U ��vZ�O�<bK.����72�(ko7nGv����E_ob��f �si�xC!�G��ê�,��o��X��.#\c߱2�)6d���C_����Y��GΓߚL�Y#]h���&E ~��J�=�[�q�]�I��wt�	�dkzA ?�.�qA�mp���t ���4.�a�P���ᇦ6���'R��y�%��>	U�͠�5w<�7R�� ~]b��s�T�~\�/�)-$޼�9Y@c�㥅F\P���M�!����I��K(�sh�y9�3
�Sr�s`��#�g�WB��1i���.�
:&ak�~��Ip�+'��ǔ����e	t@-��o���R��%̺^�Y:��������Vș;��<�I#�I_���"aݸ�����Tя�Ύ x�u[{�̾l^O�*X���`~'��7 �@���7����;7���$�:���%����an� k�#�v�L��9Z��!� UdN��ֺ�#-���u(������g8{[/t÷~�/���KE�/��(���n(�|��v�;��Ǡ�Jz�] ��sNi��y������q�8A�5X%�Fr�u�Ŗ_"^lK�%�U���m��@�+h�� uiD �5^Z��3Ԗ����2i�OfT��FȤ���^i��c��?|[#���o/�6b���co�
E����y�o"^+Ap��h9���}����?�HS�Yۈۻ��&u��|H9��g����β�9���Gi�D�&�0Y�Z3�!�[��W�����\a���'%�ָ/PA�دY��2��"�D��������������-@?�(�uUE���nH���>@n\X,6L}��N>)��]�534���F�t�l# 3y�_}[@�T7߬fs�給���G�2>�����v؜���3t�D��eM���S.�C ��&���#�� CSu9�Q�]bΩ{a�����C!1�.�*6�C�
��K�,��1�uX
�D�o毦숫v�d�'l_JY�)��gt}(�L�A�l����W�Na�G�K�P�'�#ֲ n��I��B�����<�͏��b��j&��ـ7uW�El�Db4�b�.��y�^'�ؗA�ڦ''�}�I44���#�P�: ������X�kÊ��`�a���?�M�`�|�
J��&�H�HjҸ�'�|�wv�F'�߅����9�V12������5��{8$�SM-&�_؎���� b�h`��y0�u�7e�7ޔ0�;{��W����]?(هV{�bY��t����Z���ǃb;�ǩ�Ӭ�X0k�ϲz�G�.��r��hd�>�cɲܚ C�m�i�EցK.vU�����~LT�����c��X�Վe�T+�d��Ki{�i�+k���$!vF��2n}����;��ī���B��0�ۥ^������F�g�sq��Ԝ�����R��� XN������D���b�)I�0 �����]�'�h�-�o�%!�r	�Z�w�w�!KS�����
)����E�V �9�3ϑ#=�@c��$��^؍k�ؚ�"��1@)���zȣԛ[���3�N^s��Z�È>����%5TO!��iF1j���U�AYPu�&Π)p`2OZ�b%��My�H��O�Zl��Q�l��vDpe?��Ď�k��݇bC�|y������*��Իꤚ��"�_;[s�}L�>d�dֈ�=��1�SXjC[
����UUb�y���e	��۾�l�h�lvV��H�FL�+.Q�������]N�V���J*���[
�5��\��wH�w�l_�����p\]��N�M6�d�4J�M�Ҋ�����tw>L��k�lǌ#�%6+��ֶ�Te\{���K���-�9��~���#ֿ��^�n�#�(���<~��Ev�l��>]�,��r�v��ٱ���U�D��UL��Oc��$��JJ���r�ߚ�9��x�_fe�.�`�T�$�ߓ�C�S�(�"+-�9���c����?��:��*��ϣ�4���+��y"p��8<��Td�R�aEP�����[-������oE��c�6�:����R4A�Ak^�H���κ��x�����������g퟇��_�ą��!u
�Y��r�e-�9�$�D�F�'�t�D!i��.��݉~��=�@�����~5�������ڏKݧ��q�B�lݸ��n��Ʊ��;�;�<�ıj%1ŀ���s@w��\�Xl��DI�E����u�a�n�z;&��qg)�vb��#�G�<P���-����7���1}-l�ȟB�?�l�����PȖ�e�g�6���P����<�2MU�=�	�n�����fw��՞�i��-�Wv�oJt�y/��I!f[>w<��3�8����F�p<�ks�v bQ�̻|��n��w�6�Cmh� ��ǰ?;7Q�8��E��˛:G�?db��pߦeG�&�)]�{-M�;[�S�g֮�Uk<3	�P)�e��H�F����"Gw�������C���m��e���Ѫ�*�� �d6l���[��n�����toW�^�(�C��щ�p  ���W��.��E�ҙޣ0(lָo�kl���1���0tiu�Mte�8�^궮W8����d��πVfr4m���9��L͕���\b1�r;���+xؽ�;{g���Bh�YU��B{Y��$}5؃���Wz���Z,=��T�ުcp�bi��q#��M �hV��v�#x�d�4�B���6wt�~�ͽ��(�E��+y� �{������UT�I�+�
�w��7�:/��,E�u�H�����Z5%i4��W
�mt��hn�O�:��þ(�1�d^�|�:ʴ��\��6N�ġHn��9���J$�� ���J��(=``�oK�ln��%�$�	���Ɲ{���up����.�OT4)'#�:Tbm��H�^q� |R4�[�[�{���O����ݶXp��@7%-��e�kŒ�%V�;2�kS�JG��~����F	�-8�ַGϊc&�l���O�] �]�1�*l��N���+�Q�-�[@e�(hG8�y�S��r�"��Q�(Ů�[I���8����Ɋ�s��ތ=+�a���(�!0�N�H+���&hC�I���oW^?�.Zs@$	�*�׹z�{�h�Å
��ZU9�z@2{#�	46yi���__����0�_-�Ɣ��������1yu{)�yA��r�2|	��n��iE��)���?(Z��}��?�9�!4z.tu�c�j�~�-y�*I.7��e���ӽY�*xq��������'3�O8l����E�k��v��Ƨ��F�#�("^`Uxv�#�w~s��ׯ̚��L��G{��m��t���Хͫ9t�{d&����s��R&�ڼ{��m��a@ew~C��9&�[7K-n�@^5I�j����WBƙ jvצ��&���SCYj�pv4t����(m����rd�_�%F�=V���/Q����7���>y�ߺ*�l{ÒtQ�V�g���F��UP]����5G�9�Qa���&1$<I���ә��;�����െ% ���̓M�`��e)��2K��>us�k��./�<r�-���̺jb����H���	����$/�)����y��`�7���'�Q�~�M�o�����G�N�7Uə�vB�����xsN7�\���j��Z�V���'v�>e�@d&f0�ƌ!� �
l��*�M��Nf�K��<_��ؘ�7�� [e���9������� y����rG�,`�Cn/�q�͗ޛ�Q��&��Q�ָx�
����X�HV�i~��B�lu����0����W�=:���^���Ֆ�׳SCxZ�o f/݋��?��|O���H��go\+4�~`�%��8RX��	�,���$%%e���"�t`�A��L�^n��l�����]̶	�C���9�;@�P�O�W���� h~2Ԫ�DL����XK�?h�j�1�FXe0��j��jy߱qLE�3Q���Ioj�{-^��{qv:���b}4:���E�kLg҅<��Rؔ!L��w �|Q/�������Y�e���5��fK�̳�c�{�W]ے������Og�����NN-�+�:��l�Z��ow����|�,9Ӷ�\�ä�qH�+"��N�}��J*=��V�/b�n�fV��3�R�[��֚�Gi:{��G���K�Ǜ|l{m����$�)5w��z'���g��\>��/^��Z� ���.�v��������4�QT�j����~"�s�'&�h��o%⪁�@�Vj��YZׅ)�v�a�����Fm!j��x�eq���NPd�|�����g���~ش�Μ
/����ߜ���C�s�%��:ӊ�͡�t<�R3Z�H�̗R�Ď�b+1N,�.�D ���@CHn��S2�*ڑ�1�u)�a(���4�[�]M��[�R�4.0�KvZ�?���v4�y�5�{��-.V
`��O�;�kKޏ��]
aܜ>��E��il��H��̫�Ο�3�(0,�+��C���U(Q��sZ�\�N�u����\"��ǘJ�O��oq�]��]Bx|�茏�/Uj����l-vt1��������|�������]��9��7���ё�l}�'�c��u��	��{N��������,��<52�4��ٞ:�1���e�V��|:r��µ�D�lۨ ��4~�Z�p�e@l>^4�"P�Ի��ȃ�|)2'*1@�$��u���*|�"��y�h(,� ���H�N�I��ep0��D��� �t��cI�E���	�E����� }��;o&����U$���P[
i<B��k+�▀&F��`����!�����ǅߴ��fc.��@l�-������Y5��p�l/7*Ǖ�,s+�"	��_W�t������}v�0ص)��V������Z�A�z�����1B%Gy�'y�8���5�F�� �}^5���U;>Y����M������Ѓ[��ȹMO��XG�8冏���)\)�R(�i�cG���(+g��V��/H�F�¬O�FX2ߏ��bGdb�� �x���\������݈���r��oXX4~Ct1��n��hE��#"<^�4N#��9q�d�X�S�U�5朅_�u�	�ˑDJ3��m��\������w��%���4}1���$Ȓ�Ïo�80&���L-��f��w���G�	��F��[�Um?CY����n��_j�M"����%	���m�f&m�{�=$��������@�NM�{CW������լ)y��A�5]7H)Y[��f��c���f��B@�`5z��QX`$�y5͟*��S���c�7���4�8��� �kʞ�(�V����B,�Y@eŒҞCOn�8:�g]H!N'
6@#�6d2=�9`p�	Z��k��Zq�p:*����2E0�f8t�e�ؓ[��6ׯ /{�TD�o���X[wTM�g2e.�v6:2��O�����"?����������9|�����c�A�=��0�\���P=�,�����0s�����f���] �ɼ턾�r��8�̼�g~��s��F U�T��&E&'�T2���}x����N(��_�|�~֋M
����J�Vץ$c� k�ŢS��˞���j������[>O�5KA:��d��PHK�3Nk�c[(8�2$ő��<5�vՃNe5��{��s\��usp��VTy|�鑯���<ei���<�������O��{�.d ��Rum�Z� �~����U�LLQ��Nԑ[�)���M9Sa��e�<��̹&x2�����Nʼ����܊	uz�C�?��͖pO��}�k���^�5c3����cP�2_�X�xȣ���ǞJa�s����,)7=J*�� m�Fܠdm�P.�Vu�;��󤲢צ|�k|���.���`Gx:%� :�r~���6[�y�����Ų�|��"��0oŒ{���o,�u.{43�J�#�]���ɼW=�m��`
�9��� &	�[�}'C�0����ؿ�+�Q��)VVL\2����z�aH�߸���n�OUnF�'���I�� �-wJ+��
8`�nM�Cz�,E����We��S��/�ى��{AX9�o]���Q���(�����^S~,Գ7���A ,ԃ�Q<������%���U�]	uv��<�~ �/�.�9 ���cr��B�:�8;Qm�ߪ��q�������,ۃ&^��i���H��*q�Ydb��#����P�ί@�2a�Bt*��Zgd��}�N�+m�M,^���q{k�?�!���3!)}ww����1]��/��೧��b�V�W��l��;�`���sಡW�w�Z�9F�T�k��c�������UB-ά����ݜO�B y��J��B�N/c	"����)��䤧��R��6��9�u��-(aOR��ǌ���_g0�F,���s���q٢��
?�cAqn��(��G�af�~��q�](��q"uF^�s��1>T9����?;�	������du������z� ����������i�b�w80�O���w;b��P��6�?RTrA ɉ�R�ϗ�sJ�5�)M& ^]K��[�7�gn* �����]�#�'i2Z�A����  N��~��T���tE����Y歄�f[�頷��Jr���K.1�,�Ň��_WW�?{O�@X*琿q�����!���~��,r�����jn���:t��oOF��2�2^9K1�GF�74%_���S�?��hRm�D��K�A���c�<[��i��6wW4n�n�0�U�6����mh��s���=�����0�r��ԅg�ñ�HU�o�3JS.�y�3hbS��h�d�dF�sg ���ڥj+�ѝ�VAw%)Q�S�!�ũV_�o�ZQ�U�� 8�d@��G�b-"�E���+��Z ������/�yȠ=�|��	1�gz��Mt��h�gk�z�e�xzdPq���'iV�n>�`�-h�A�p`�#Me0�6�� ��p�x��m@1�Ti<��1�;��"�2uVB1@$����ƪ�|�z(<�4�&�\�&��AEi_��FZ���mfNYA
����K߿��K3�i?)��L����2�t��Ӑ���1�/�_������u�P(�l�z@���X߆�t�1���;� B-\#����䀣�0?b<��`q����\�ˁk�s5��%]V���� j��&�>c�z�2@��K6��Z?�r�䥬��`f������R%�K��L`� ��UE��v�+� |�;�񂟬�ߠ�[��鍚^�(޺�|P�ư�(�0,��I{"$D��9�<^#���mq�A�U��j0�6D���~��p|y��2�v����􋩙�U%��T���Ћ�0����Pp���|�6��c�y����r�x>W�l;e�/��M�S͖3�:n��b���+���W�j��^�?�B�Ѭ��&�TMɭ>r(���g��6�?У"_?��z��`���L�Ɋ�����쌒�㗢����z1�kRM����I�v���>��)=PuԦc�6b\�؈ro66���(a�B����V�o���ƯJ�I�u������v�8�[��<����������V(���! Y[�$����X��W��|�?����Ճ���Ѽ�n��i�����p�_����N7�}xۻ�����=ܢ�P麹�ǝ��NQ��>!}\��ry=�7��(=�[�z.�@S�tn+�beU�s�ڨ0�C���N@�hŦ'N.t��ח��d-
��'Yn)������$����a���SZ�=:���B$j�9��lEh�j���႖I�֊�*33l��,�c`��N|�����:O�����Oi1d�(�hCo��c��޻��ؿ�ˁ��[�~�T�ͺ0sC��~�M}���qj[!�%�<����&[��.Bd=�^�t /	�T�<t<UD#�s�DR��U	bxI�vE��1-�)L�`��v�d$�3z����7Y��46���{���(�CfV	��fnQ�I!�!�Y�^
�=����.J�>
��<�Iƥ[�A&9`�;֓S4�ap�f(<���G�_�uy��2"Ϡbn�ȲDi@�.c�r�BEhXp�R��\�R��"# s4~i#���Ѹqe��k 9���%͈q���+��zA���='|��W$��E�.�#G߱� r'��
q�e!�X��		7b������Re�U�F�?	'4���*�}n���j�oB-��R�!|���g�>Gܼ��	äG#�3�i���ԥ���̲�9O��եD�ߕV� ���&��El�dx	�n�2$���*x���_��0i�L��&���9O8Q �ĩ'�~ Cg�B����ܩS�ֶ��AEߴV�!�G��"���.:{Ճe������Xqog��ŝW��E���Rry�&\錌"�l���S]b�������,�xOT�����ԕ|@�_\
��^t�t�=�fk&��3s���i&hB~'�H�Y���[2]oPDL=��Z�il��"�V�J���,Z�Y\$RкĶ���CO�A����S�oUvBw������o1�&{8��}���J�4�0�.��l#�RX::bK�g�Fg��79{�Y���1�g����U;{�y<{����i�B�㑓������SW�4�0������.��}��f�n��va�LyJ6�)+��*"��.k\'�tj&�&��._�������D�嗀l��In�ұ3�o�&��͜�{��l@���g,A_r�(�A��o�)${�o���>&-��e�|Ŗ>KhΑ�8if}�$<.��S^��&zC.HC�(�(���B �5���;m�ji[�c��)�x���[8��~�������=.N%ja�.,)�,/�U��
C6�2�=�Ȃc�7A+�*�W��L<�L?NR��!�c�'��p�{��䟌�_��@J��i��gځ�&C��S]��M�o����=C8Av`� +����;�
��b����پ$SV�*�O@�Q��E�A>�*@����[Bf�b��arB�[CD7���ū8�v��۞3��&��\n��z�s���|x�����
F�8A`K�[
m� �֟K��޵y>�&�ҳ�|�Y�Rөsh��L�����A��Q"Ln�-S1�b�e'M�q2�����w��~��u)́���`�/��X��+����Nw��Đ�C�"m����"���[������GrcꡌG�߶2�ރ��[�\�u]I�_�;�u���̑H����Hg��@E�ޮ�M��#�SB������z3����֓����-�F�a�P�b3����d�=G�/b�>��ǉv�����U5ԍI�ޡ�A��a-�޽3�
�aࠀ%؄ɍ����'r�,�i_�h��FTX��R=�D��S8�0��_��&�Ыph�a�h�+��3_��P
�%����th:�����y���[�YP@��;�=�������>/Tp��ҳ��x��J�2S��ɶ%�NJ s>۴%t���hܼpe֞"QY��*a�vR�?{9��&��2��멜b�bg7S!�3Z�bw:3<z��`���q%�=��A��]�H.\#H�v�G� �"e�(�g�,�n�GG����[�	�7X_A�x5@N���b�RD�X�+V�[I�!�e-��\.��3�~�Z��
�ǃ��g�u7�RV�d4,"+��1������m	��k�&�0*��י&�Tv��ˍb����"b0����|�xW2��rR&��W")�W�AS��F�	0n������ߎh��+��y��џ3C�>�D����sm5�k���Z��^oEg�E�r���l¨c��l%�>ψ:`�w:��� ��
��9���N��˦&ǵ�����^e���4ٯD[�;��1'����C���S�\�(�F'G�@-M�HB5p+؜O�����ՊA� �S��K�>�D<A)�~�U��(�\�8F��[n����{�r�[��k��S�<�p�	"?�r@�H���ɚ���4!�����Z�K���?���߹((�(����%���8�1��@����ԓ������0b�7���l�wZ6������|��!1�į�$2����*��֊g��T'�Ȅ�����Oj�>�i�(�\���p�_�\炊�
�j $��E�-�d��Gvq���xCp$���bGE�ɨvŐK�O^����~��0Α)����Р��;�J�(r�*z�Q�G��A}�,�sU�5�kw,O��?���)��H�fϞ�p���t�Z�<H}ʱ��%��ꥧ}'���%U/z�BF����3A���i��+Hp{�t�T/κ
��NG�N���o�ޚ�9{�������G��~�<~(L�Ca�d�R��(@+��1�߃m]2���&q�}�F�!��v��:�5u[���L:a&���N��hx	�q��N�X�K��0;��Kp,,u��EX\f�sل��O�w�H6\b_����A����\d|^s���};�R(�7�<�i}��ܚ^�$륾��ͪGu;��#\c&�-��7��lܖ88��O�b��	a�)�g��5��B�]���k����	&7�X�w3d��g�T��ۂ'9����?�UE3$�b$u�h�E^�9ʹ����
�lҬ�j���K�M����v�'Ò��9'����c�����G �X�y/����e�~����6����\�o��9�pg�,j0�������G�r+X@�#���o%�F�\������n�����Fo2�����p��� ���R=��,�&1<��g�b2��� ω47����l!����7p�[4�r�l��9X�E5cs��M=��z6^���nf�9�ٻ_d�Gg*Fz�{kr:����udG%��P���������x �2m�
"�R�lvqF>B������nD����5���[j�,���E���4*��B S�U�k'����mvQ�u�Ǟ���2@v�K�����q�0�YJ��"�P��fo��E�;��ӈ#jCp�F�J������w/)��J���}��H���T���-�%U<�NLv�4(͐���Qq �r7�0I�)�R@i˲q��y*����H�͈�4��l��9�[e��s��V1f#�L��>��^N��a�?|o3 D�l����2u�u%���Ӿ_��L�ڧ�H��糹�Ia�A���@~��u*D��W��5�8��}��V�K��!!�0�	�Ӑg�˦��O��_񸮉���pS�p�Y��ӈV�h^f�D�jșo��e+#t�Ĩ+�8g��U�B��>��IS�w`!��q؆�1�|��8�ӃQ_:������,��i���-�l��	���=��t���״���Qa�Â�+��r	H:�T���!�͢���r8��ˊ7�^�c�C� �����H��Ԣ�L����
�yǦ@ ��&K�b_���u��2研
����Na����7�3"1I�m�lua��8��NqL"�P��@^�Etg�J�=yC�BÅ�>�c��l@;y lԵ�՛�8��(!6-�fm_$���&`���7X�&�q<T��/�$|��V��^g��2��'=n+����ũڱjZ�㬉��� �}�m�'�!�STFdf�:r�~���S���{��j��/@e���Mɽ92 ��^��@�C��l�_(U���=U��Z�wF	F~ ����@�0�q�x"����8��1�j�ڟ���'?
p�jo��1?�>�WZ2#	��K��QBe�.��{�u*�>�\ئ�Ź�Y.��������?�]�!hwS��&�3�EK2��SV��iH	�=zE�G��s�G o���3����aOD!�X>p��4�c4b�?�w�^�UC�� �^R�N��닙���e�H�����s�q�K� �=P�����5��W7��lipv%I� �5�'�8�Ԏ��������Fm*�UIxp�h�N�=G�\�%�|����}�'��,t��eC�!��ӭ�z�@�@V���h��|AaXP�^�S�W������'�Mľ ��H��"@�|�㧄J���B>ji��=�fBh���~��"�8kU����=�pk^xs�qc-'��_�j|4���0���u$ߐ(��cːF8����ΐ�1 �V�����"֕�,��2�)�h�����{�	;�ի��BT�����&���r��~�S'K7*�c���(��F2mL�	�;�� o�9t(t᩵����G�<�g[_�ܭߥ��!+2��ұD�q4�_Wai�E����6������1a��`;[�&�I7^~%E��f����f�U? �y��6�	ރ��\�b��=)��sEw�`���\�v��
��|sPؠ 'C�����?ݖ�_���d����G�w'���>g���`������#L�����|PZ����)��lH��v=*�Dxཟ�<�Q�p��/)gs����YZ�M��ku�(�����>"��6Q��\4h��,�d"��H�K�؆NRa��F���`q����cu��(,S�߾f�w#��rp;��oCF,��gi�7���c�$u)Ys�(�%<I�f\6���h���}��p@��l>�Q�ϼ6=�E�s� �-�RV]^]�W��%�O.�Ż��� M�wZjA�o�GP����~Hz�&|?����\2�������@�`ߎʜUv~܅=�L��+S7lL{� ��+�ǣ]��6u�׻��?A�,n����lͺ�M��=�`	I���en�_aU�Cd�����EHj�#�.ȭ�]��PK�\�1"�9��a�v\o�S��L5��ڹ�J���C����V���Ic����nG�y�|7\Ͽ���=�l�����c䢔D�rE������(��k7Y�� tT�1��V��(��P�2E{�� ��J(ͱ��L�f�fq��Y�(�'�P�g���ף��Zo�≌`��)_�e���k��� ���d\�Bpŗ��j�X��";���4Ʒ+7\o"�$�I)¨L��L�.� �JC`W�j����d�"�,�Qx��?H����հor���t�3����d��2頏���Z����?�_���@��N�p�w�c�pd�����e��Kݻ���9�@J�+�,��l���^�g��:%��DBF��l�������[�j��h��3e��͡%�W�χE3�-ܿ+=��(r�׫��wa8�#��w抺�?�T��
�RP��JC٧J��(޼�~q��c_��Sk��[�f\;��wP�P��,c?��?�@|6���.��)5H�I@7�j}�{OGI
�ף��������dR��&�J���͘��1ocDϟ��G�$&h*]HMߤsBas~�e�`$�~��w��++ӆ��5���2@�=���3�����)��-�7Y�ά�@j��� �H<��4��N3d�*j�0�IR���I�|��^��P �"��@x�w%��K)�A�e��Hg~E\���y/�Q���GL��׌�����~��\ע��m�8�ہ�}�@�c����|]��#39���6Qc�CerKJ�-nk.��UV<���J��Չz�UWy��V�{�NCﯕo�R��$�lOlh�7�N��W�ɰ��s?H���S1X7�Q��앆�;��F�[3��c��kl�e��_�*g����P�h�x���D�t�	�_{��e�fe�g��v�*�Dg���O_x�����G��C��,ʇD��B��-���@Aj�x\j{Ԙӏ��~.����b(�گK�	W�Q~�����>O�.�N����YL��L ��x*H���<f�S$r:rB�I�+L�@'0���׀��r�tʢ}��"O�&�O�Y:�K�
7=��/W������d�����n����p/�:���,���9r���L�d��^sJu~x�c��0y!w%z0�1�ٮ`"&1n��t�)y:��WR�ᄣ��J���hy�Kn��#ۄ�E�2��YS:��R�ݪ��R��y��^�z\R~�?�{��Q��,�;����G�����}4ڡ�B�X"ߙ��Wڝ�=�Ș���DḘǿ������B�-���D7-3��2�_Xz��O�${8��������[�Sc#w��k�$���jj!�,:N����Z�溝͕U�]��,���w�����"4V~̫�t��P|� ڱV���,`m�z��>����?l�(P��!�#��F��-���N$ghE �8��w��Ѕ̷����ِ��<ywQBuu�q������ɉ��0�����ts�X�+�G��؃�ӋY_������^�E�����T@�r+bĺG�j�RP �����󡈧��PQy�a�������}RZ����H��j6�	Q��3q���Eӽ�Y����?�{a�5���¶b��E�,�%�'�>Ó�����)�D�����)v�g�o���=罹L�[ǳ1�`��-��˝����;���,ǲ��PLz�K�M��`�ѷ��d'}&5u}�����q��s�$��ROi�@�:
:=gh�%����8][.�P��4H^ *C�ރ򉬢��6����4*����~s�2��P������z��m3��[b��l{o"T+�*�R��3��R�If����8�Ytb����Q��<�s�����~z�4 �<:��T;K��9�^0��??�����Q0O5��OR-̊����EEr��=";X�2_,^�D�a��6nj=��`6a���D�3��P�2�� ��Yi�C�!C�M�)k�Qc���3��r�]1 ��'�9������j7/�RdP4�H}%�%o���YZ�e�>�0�$���;E�H7^���~�AXz;!)����0.X(��;��w4���O&T�o'Ǐ4����.�3��9{&�p���������a���k���N�1��P�����MoP��
Oƃ6�^>�I�<����o�:onp|b����z�O��6������QZ8K�|�vv�h@a*�co��K���^R�M=�
��fJ�<U���j��*�_坵�A�y�
��:7��I� �Bk&cƵ��?�J�1�Y8���A�+���>N+��эʴ|�O6�V�^�/���Nr�r8��b�����Əq�ޞ�i(�S^b�5�#Bs�Y���++��\��p=���>���uGn��Y#_��].�d �����yI(��"l-f�}����-��
�+%?�����{T�i�a^�A^0�\�8�(	��oP���vLv��l���_���j��\�$���q��F�O ��d���xf�&��F�q�Ee�e\2PZX�2g�����SCz39ۻ<5{�$����t��m��4����kA�-�O]�ı��H���
�m�܆:��i|�~��Ǎ�T��*���ԅ�[ ��2c�+e/̦�z3R����2Onۿ�Շ<]ppD�l�m�o�A�9�4��0��.G/Q�#|���g1�q��CJG|�J�ˣb9�%g��`9�Aݫ���^�D�0c⫉	�{M�.�v�%+�7p~���O���|6��I�JaEqC�*#a�R�������w9��W4��3'J/��>��9�/'K��n �O ����'u��C��sʦ�0.^
?ij��%��ڎ���A����������D�]�����q����;�|^�Z���˟b�hMz�.�Dˬ�6���BZH�]npn&⧤"g�*�=�u�]�d������\����Hc"�:3^ �7Z5�g;z\��B��$ϐ���R��9� `F4S^8:-C�ҷ1���yt��Rs�������`~W_�]�$���f��^����c
��֤@V�I�|��v�h�)b��p�O.Z`��f"�>�F{�������$������b���֪��D-a���f���\��-���\��J�3�w�����y�2��y8d��Jq�!|�-�i����2zf�� ��� ^���Q|�x�)5�Ĺ_�Q�bV��0\v���&-zFX�p�v��Rd�)�ttg![df���b4�bݞ���b[k�E�3];�N��}-:�A^];��I_�U��_���氻��S���,[ٽ�0����[����"�J�>�H�i����SJ��.f�Ks����3��v?��I���E85IH���rg�O�'.l^�O��q	�YCU!v��+ҁ/�DRRv���E�!�T;�X�ã$s�|�*D�M��X��r�TАdr`��"R�Kɔ�N�U�`e�����F���h��V�}�c��!�:��S��W�7�	�!-T+�zE�g�������!��Ϻև�-�;�c�7;M ��5���I�"@���s}�=��4���c	��?��N:SQ7�֦�b��]k�����H��g�58u��W�i�"�m��vF��,zC���i4!z����dG��r��`��V�syT(7���I�7��ALv���r���|��]\���IK0w��gI��v��G㭑͡�2�Gr����L��8��e� �����ٮ7��]�G�]�HG���Fy��B���	�8睳�F�w�s�[�Z!���"��ԅ�?�cI>��W�#�(0Pz�4��oI0!�C�
|��k�}Fz�1�j�N��<<o����ݴ����Ƌ�P�$;�%�Xz��B�.�+gC���_'LD���O���$e�%6c,�g�`A�1,̩,b�b٘���"�9��0���A-N��fc�����{ǈ����8J��:l::��X� �a`>h����<2/.��ph�	8!�4�����ʴ#�5cєsU�j�zý�V�?_���f	���A��+օCn)��{�աA �o��ʶ�7ׁ�S���{޹�\l���WBX�Sb�OsљfA����|z<uc�H^s�IO�#�T�<"��J�Dx�쨆�H�md�y��k��Yi� ���XYn����VaN �I��D&��w�.�&t�[1��ǋ��^Ƈ���W�g�E��P1Lx��03�JG���˩p��s�&�N���pȓGg��<g�����6E�2�?�F��''�A����B����F��וd�v�s��t1jA�J{��z��F�����3����#��q�`��f���K��� ���	���{m���]Ri�I��C��j�}C=H˛����Mq'��(���K�����YK4}�R���/�Oaz���9��=K���l�h00���P�/���ܢ�� ���yG�qk��S�J�$�7[�a�@��A�s�}��v��k��O��O带+n�8H
�x���y�~�|�S���I�*me�eLy���\���}H�����c�H��1\d�Y��� ���	s��^:\����J���"宬h�c	�e���|����1{��BVN{��Iۜv�r~�Aԭ�("=��e!I�|_����(�B�����=�{�=/-�x�7G�����z�v���x�޷J�*fDx��٠"�^��4=�D����xv%�Y"�:0~���䌮�&,Y�?�eT�u(I�81f_�,�QQ�����Q̩����]!�W��ǀ8�Z��1I|bӦ���[F��a�A���=kC��Z�eEt&ծٞ�Vr������S�"��� A���+�����:T�v3���>.��߫=F��0¡��q��Q����)�yO���y(&i��KY��,BD�QG���z��"9(za:��bZ�r	��Ů�����+p�nj���26�o	��8�r�
���9of�)�~ �Tc�N�'.l�{Ń�d���x��L���`:&P��~�]��O�cց��@Gnr�x1���1�]��t���{�xۘ��d�Ċ�k�D�s�����f6p1�9�,V��2cck��.�R`i�z��P���6��
q7���yB��vO���p��\�m�>�)��$$y��� �h]�Z!����@6U�+�K
�2��&h:=��eyu���k�w�.�j"dX�.�'�a����O.Bb`6�~�|�/;huޱuP}����E����I���!�j�#`y�=<b��r�h�d�cZ��mΜ`Cd�#�a��ׄ`8@�4k��L;�x]�����C�ɠ��o@�.�A�����b6y�bq�Da�'�U�p��Feo����x"�|��Ui'����M�c(��[�}�N�h�����7��3݋���x�V<
���ƈ�4�ƃi<���:v���$
<����5_�����F�֗~4��]j�lz<t8��/�=5ȸ��3�2M0,�8������=<}���$���'�T�Wٓf�!r���(x�gj�p0%݆�Ak��9~"�٦!�&F�o���w���PWe]��wer�&��ͬTNJ#u�|�!ۂ�p���$`3m��9��q�����@�2 >-�������/��
��ZDk���6�@8��#��#����'f�����8�č��f��:֭�k"�e��O�%ˋ�e���������0�$�{�iV&V���?��x�������g�����x�0�?mi���[Hl�}n�^�8�o[͡�}ŗ�GW�)�Q�zc{�%`�s� 19�|j���kIƻ�h|�!�cJ��(��?�:W��ӵ�`�X#��a4����n�Ղ�̾�E��� k) ���#ԕ�T̮]�֪�3�LN/�hEC6~�g9{��P[S�``ªg&Tɗ�h�f�H>�x�����8���I��	����S_�/�{ ����U��k<�[����6����$Y�Ϛf�c�a�27�(3�)��5�ʤ���v�������P�N;����w����ي��D� )~��fb2��%�W�Zg��,�Q�'$�Z����OGp��h�!��i�$nX�\1��G�;�MGfǱ7�����\)�D-�7{2:���m��WJh�׀j6L(.�O��g3�� ��tYD$6g<;�w�N��:+��7S�9(x�Տ�62�hXt�`���jxBϜ�y�GbK�������ˉ�`�<siZ�!���W��X.�OR���|(h2�H�ӱoV9���xS_8���]f���KZ���,
MO̘\۟�a��Ma/��E#������$�ӌ=���qJ0s�p�6 �Q9����G�-)�)P7�1F͘�������lԣ��u���(���C! Ǚ��-�A!��b
)D�_̰�D��\,�;�p�U_4��R��|�VF�~i�)�v�+�>�\1�0+`/�*�Sr��*���%���9�ل���[آ�/]�rnnK��X�C.�3������ns���h�;�;9�ܴ��� 9+O�9�B��+MC��E��Gǝ��O�I�g��.��	��G�MUN�}��1���B�2-���Ȕ�߫}$��m�F���s�|���(Q��;vb��H:���Q.�DQ�dD�Y*}�d��`^���Y����6�헶��A����� ��%6!��*OE���_5l����)�B�іE�������B�����5�b�ϙ:t�_�(J�Ҳ�����_�OR����]*D�� ��L�X�7�\o9��V�*#�'1C#�"A_�����Ҝ��_�@�m��ul����eY�O.��K�����*�� Q_�$�2.�9�En���P��kԧ�o�ӺXQ	�*�G7����[�b��P^B��]���ק7�����[R�ϲ,,˷��$��7a���t�~X���Z��}��T�)��d���,�
���]ۛ �;!���Џ2|b�O"����ǂ2��e�z_I
ob�3�}N�&'�;*����\��,��yr�����'�Ldk�`���NxԈ���x�V0u���C�Zu�(�ͨH��Cyje`�hǶ�6�ð">x����@��kH��Ŵ�E�q�p�x�F��x+ч��y�#�n��\*��Z�WR���O�7�E�T�f]wo�pX�R1O[Q���J#��~c���|N�e���b+�A���w`�+�j��ե
_� >�cZǶ�j�3���6~ea������;id���&�Ð���z.��ЭZ�WAh�84-by��ц$�_�j������ؽ/Y=.�+��~0_k0��1Ƣ�s�.�AKC�9t1*r�c�<_��Lc�}(�G�����D���H�S�I²=���q�f�BE7�6F!796V�Q8���h�7O}W��d�����|o��D�����|Ǥ>w����$��������T�O~��¡",4����Ks�U�۹�f@��o�r�0�c���w��3�P;�S:��K`Ф߲��^�))9��DdD!��x��6�������3�jG6���YIA�L����T
=+~�߸�(a� �.K�����37�:����W��l˭/ؤ�i�@��P��Ƽ��k��ˮ^Rx�m��=FO��U��h�����7Q�J�o��#t�AB�&Թ�x�}d��վz">�az�����[J�h��'�]�P������G�Y�X�Ҷ�� A&=��d @_�$��5|NӞH���� �{g0\Xqмe��򴢰CP���G��+J�=}�T�i��ȣ־%}��Ђl����ݟ����
c�*+@�P�*� Y�}@ �'%�&O�WP�A����m�5�Rv��X�:H�?�v?�/v��ػЙ�RJ�
��S����+��вDD�U�>�(�D+}���%�Ft1x�CO#�[|��Y���蜛�%��wD-;�2�z��Z�e'����~���'���6���ì�����7�=��^8�C�������F}�&�Q��{鱌^s%�Uex�`��J�����%O^P�g*�ae��9oى��b�������Bq�����`@vC⢿E$8�&س꺪��`.}@Ʈ'V��ΰ�� �����*�c��� ��4 �;�7��g���<`N�䭈���k��,�`Á��a�Y�Q����Pɜi�}��<
i*����&���[A��3��rV�B��,�N=d`d0m���ډ�q���g��v����1W
������I*�����eÃ.S�B-�a��ݹ�����{�Ea��b�o�R{ǒ�c��OFNq!�l�aҨ�g�9$�"�ˁx�S��/���P7��"�6��1���kF�KkXhwxjx��@Dǐ󱀽7�-�7H�py�%��MP�cI�t�2U0��g��)���qή�@ �q�f�W�g�0��(!�&A�+Qt����?/���"�3a|��GVv$������&��=®-����cI�ͦ����7L���9�G	m��C�v6��_ou��wV��d�AAk�}�d4�X�ɚN2����?����	��5Ww��y���� (����"�` ���<�t�g���&�y��;��k�%+R#sKi/9����52r�co��T5w����L�Ex_r�RE���{���R�IT̆���M�"�U5�sF���2����}�Q�X'��w��A�\p�M���¥��4xD�9?q�bS/9
�E	�{�@���5�a���ۜ��V�w�6�p���)�ޯ�R�e�!��36R[����Z'�B!���	+����[�r��s36��Kʸ�USb-~��ߜ��Ӯ�	([�n���|颅���o	�m�3;{���77�Bl1��g���a41ϾSBn���6,:�6R�d��2_Nrn�Wn3�I�d��{9�aP�_�E�	�N�;����#�o���-s<�H������1�1�9H- rs������w��'�0S9��-�2����#�H�z��1fS~�X %��
�����us���-I�fVo���TU��C�ϔ�M���f��<SiΊY�Ȫ���F�j5I���ߛ��^}�&||�8�r	t��"Lo��Z���> �$	1����:����M3^/��0�^�����c<��m�T�����dX�d�V���>������@+$��j��X2����6yB��y$�;��mM V:e��pª�mʪ�����gGx�R��r�U�F��j�-���߽eW�-���\����g���d�^�!k������7�jE�DM��
�<�"�]�km�}E�ȅ�0?4�@U���G!~,���崂p]�ۈ�H��=��160hPx�o���L:��[��3�ˆ=ʚF�6:�2Z]�+�mj�hU7��I�k4�`��A�s����B�3�}��~>�;ɡC�0�n�఩���PJ�uəJjz��3o��A8b��!݃I����}�?1]�B��a#a�>[Iɐ|4nXN5�$�}�:�})���b�z5ny(NE�{~�삜����m��R�͛c�R����n�)P�9k1���WeF���KS`�j�r/����g����ܡ轾S�O���r�u��	M� ���ǑS��i�@-�N�3x��=0gHT8�DG#���)�Fdv0�%6��q������Gd9�����g�����/���O����\��3c��[�7��ri��)6�4�.�;S��d)V����Pd>�'v� �TGX)��P��Y�|��:��?̓CX�AzlF�"R礮��~,�1�,�(�^��V.��+ӣD��E�E��go��m �R�E+�)*<,NI�:�7�[j�X ~�$� ;Rk�a_Aؕ)��������XE�j+�c=<;��}5�?��8��4i�M�Ε'�Ԓ��u��I�xh�f���M���6�$�CRs�{y�tRo����}�V���M8��e'��:�ٴ�޳�~޽y;�a,�^]�A������7�POy��%§Q��b���BA/��v�a�u��,�B�|tj�[�Ƽآu\���ŷ��y���uƅ��71L�	�8��S-�����t9z]���E��т[h��/h���97�9����/bjMQ�Hx��o]ǡ�����Y/��� ^���_ Z�� ���j\�j�^��jj�_����J��w�ѧt���a��e���$��7�W��I�@�����5U�o�FߥkT�9�28H�C��A���ї,�X��V��4�u�ˏ����8jF-��T���5�vñ�N�X��)�� �&�����g�u;����7=)Tc�c�K��X_.��A�$�܃>�]o��i�\�>k����4۲����;p>�9���������H�R���"% �.���.�1���U�ׂtT�\?�;u���]~p�5�F�S�WJPW���H_1d��7��� ݬ:�@��H�@ꊽ���*� O6	�m�fژ��o�@aJ?D/I��47��\D�fD��SD��?�P:������o7�2����Bxc�ͪ���bu���ydYŭx��!}���>�ю�Ke�[k�(?�/�.2p��?!@�Q�a���1���Q;Tǳ�<W��ߙ��rf}F ���q�3�l����F�>���E��G�H�=��R!��=, `4��Ve<��Jy��*�h�Ԏ�P��<�BG߱�L���!���eGcEx@,��d�u9�CVү[Z��o���8z�ĆOeVa=��Oʚя��j�ADZ����l	P�qgV��?�6�`�
�lg�?��c��zq%
{rѨ��b5�|Ԕ�_�,����b�B�$2M+��|��c�8��t=	�,�r��>�X�%�~��S�kE?Y]f@����0T��l������@
B�W2*�L󌸣;1���^��#��&-�	�6eZ�Ή�Udk�_L���X+��NK���']��" *�T�SG���A��G����}iYr`�yI��O5��Q%I�����z��#�V��/�q��%[M�<N=��K}o�%o(�Nmk��d�(l5�"4��7{9C�|)8H��:�w�V��ʷc�T�+���0$��>}Ӏ�����EЯ���=�v�r���5�^���E��X����-N�]�{f<�����������-�<g����|qW��wّ2�%�	�6 ,/��#ۍ"�����z"˰�����k�f�AC�V�%$�*�c��{�=p�M?Z�!��r�?w�(� |�?�&[ո�)�/ur�u#�(]dZ���^_��֔Z��Yp$�|�IK��t�!�w�4���w���cB=m�.mw���g�!c\oP��\�H�������[ʸҪٍ�^b�lo��������f�v�m%�d��,# � y�br|�v{TN������U��e���q�&/J�«����/�CKy�r�vl62�����u�3	ɬ8�L?�bx5z���Ba�v�_s����z� =FXĻ�՝F��(?�;�����>��g�[Ç�t5p�)�n� 琁ݟ���vk��e?2���I��dPy�=q-��N�s�}��������D�O�[��z ?�Ȃ� &�ܠ��v
yLq��^x}��S1bL#:�Y��q��A=�'��X�L�\&g>�;F�]�W�G�;вܪ�b�<�\t����v~��_K���3; �Jnֽ�tW4�z��`�Qs��&[���z�����w�[�n�ƃ��J�m3f~|8�4J�
sY͆;:�Դ~�Q���v}µL���|��A�1���w>�鲏�����Y'��i A��[�Y�f�Y�ԡ�T��UU`�Kǳ7��F�d"��M#�\�Lz���|�Vf�*&ZѰ�T�5��A�C�\���A]^����>��,���"�Έ"����@^6���B��)�(}&"��Y��������-����(�a��N�5�lMG'�k��B��6s��ݨ��,7@E}/hN�1�ȑ�,��JJy��Ldf'�OJ3 {�G+7����I$������������(K0	�#0�y?��Rl�5e&_��ڠr�9����U��*��*���yގ�\x˙|��W6^�v0�	�"�"�ϒD����� {(\���T4���Mq�U�/��s�N�2��R>;���k%����\h�߀�!<�V�&��?A�I��R�4��?C�$���H`x��"����E�U�&����g=����6!�_u�h/.�ZJPu�Y=e@T�T����A�I�dN�h�?5�����%gY �әܹ��,F[|RR3���6e�E�-F���0�O��;�7�	�ɜc��+�m�"���O�]V���E��g��cZ�W�7k���w���e[���/?��4vLG~�mbl��3]N�FM��՞<�C�� e�*p,JJvI�2���� =�)��:V������v��K4��T櫅]��^�PlX1W�-1*Mr���������F���TZL#�Ӻ���"qC]��)��)@�'�E��}�U�N/�&�ڪ�9u�Rx�vpm\���r�ZNR�J$N�Y��OV���M(iي�)ne&���v��$��x�6��~3iƪ��R�ѐ��0O ]����DQ�K���}����^9�ѓt�� �����Ǹ�.MN�AA�<�Q�cX�P�Z��/���� LQ���	�.�{a'j�+��q���'������������z�4t<;��TIL���dj�u|��' ���H�S�I��\���/�t������ ��&�(�V.��WX[�,Й����Pס��niA����~o��O.��
�>����=�2-��´]�2�xM���O�53�j��ZQ��g��t�8ĺ�-у��]��;?��|��l�y$���$������aH�4����0���T���j{N��!�Ĥ� �\R3���@��Ĳ���f�����*�/J��(,��dt��37S0ܷ��%: zuH�����z����-9p��Dn�2��df%%�� ���$�j�{| x赗���'�V1�{�g�<�����X�CI���������&�}�T�Ŗ��N�5��m	~�_͏��V�`ڿ	J��2y�^bD�ݛ_
���tG�f��k�p1;坜�����pn��&�C��Qb�v����N��26b֠`�7,����C/��Plñp+CW�\$U�o/4�1���i1�6F���t��
��(qGk�F����zM����S/bj��(��)�X�D���Ye��D]�Ը�toMP�7�m�̢�9�aڳA�M����&���)�6���~pKY�좢�i�ȃV��
)��'��<���O񟁁�=����$V���1��3!䋆G��^����(��04+���4��)��hdH��>�9	���U��\��ztz��j�rv*�PBn�Ϯ���l�]�BW��r�B�+|�������#nL��h;�j����,M���tO�ͪ^^[�51���P�7��}!�G,j���-G��;1��w2��B���N
]@�gx� \"���_�{´�{jX��d
�j�vo�z{�mǧ�6��ؑ��e MdԾS(���Б�dR!�c���C��_P���kR�w�rm��̐$6��=������y�V���p�6�Y�N��!O�AC�p�������c�I�͎�*v[Aj�?pT6~���.A:'��!�������4��A��ʑlt��c�d +��>0�i/�Dm�ÌP���s%!�a$�]_v�W~6���>�!
Bm֝�(��U��1?�Q�����9��Dc��3=)��C�r���3&t۴ܯ,V��ו��ʚ9y�mʅ�c	��D]�&�b���B�݌r9��|!�΂;2���yjb"��Jf���H��4#�uOz٠��x�5���������y����")�A�/���x�J��OyC��7�����i�1�a�݂OnK򛋛g37S����_��p~4mn���v_���ɾ8B@-NV�(�	�� K�E%=����TW�r&�X�	K���%u��B$��M�ۚ�Kivo����E��aF�f�Ƈ��vk;!BXw��o��m��;��V_��V�1�L҇�h<W��F}%�V���)**}<��$XD=����ԕ��	z�:��<��.V(/�Fq�>vŲ_��'o�g ���4	Z�3��@��1R!��u��9=�bjy��k ���=���F:�8���V
z&}	B�,OL��]W�}�9�Z��f>��	������P4:�!�.9����Mo�a�����<#]8���3�Q���b��T�$Фro�N�ެ�h|�6-y1Q4��rF����Nل%�ۯJ@avh�$"d������v=!E���d���ŵ��ޕos(���~�q��I��>;�E�F�`��)�KKJ��R܈7�U#�}��D�s�z4�Y�k%9�p��� iw�D)qc ����y�>[v:�i���1K�/�+m�s������Vq�C;�%��<E�M����b>*���\�"��9 +%�U�,�e�D݅M��i�g�g���q��|5������@(�1*��r&��3ò�R�b�2��u�l}z��k߳�gٲ�U1������F�����-.�G��^HY�/�i��F�t��������4�n��G:��`𵙏��j�W׵��2�?�.��r�8�<������%��H�%NT$�ѓ�4�	��hG%k��x�X�yd@��[�����a���N���)�J#��:��;����hk���*������~h��u	����֖�ۜʏ��g�#��&T�Z�l��_)���湎1>�r8_*`<ѧ�P҅r���T��q���:*E�T��d��D����C�ۻ�^�}�K�7[���Џ�-T����:R�. K�TL�WÑ�%'���I���>_�� �U�m����}��"�f�yoˬ3S�)z�w�����h22�j��˒��F2�]m��%!W�o�;Zc�����_��Dd�3�rf6��H}��2�Ro`����U��'ց���&0��*-�Um�jg�ףwU�f�:ui8X����}���u@q���L�p��T�mm��ayΓ\�rc�DF}�ḍ�L$>F-���.�m��)_G��"��b�
��-�U/1���3+Y�iTSGc�����}!��8��-�FK?Z'�+��x6Mk;�[��8 ��RwGeA�!Q-���M�aJ`C��M�}p�-��q;��+��ݯ'G���2
¯u��^��-пx���mM9F�S�������sN7e�˶�ƲǳK.�|�]0T�c>2�Il[�vh�RA�L���Ǚ�(b9���9aZ)3�.�Y I>zWOS�YΔ}V��6_jf�a�?_��������q'K����)�ɕ�C���լ�H�r�ddC�=�͵��-�j�Uu{&)�Ѫܧ�f��f{�}�Fz��1��(�z��Z����_1(Ã�6���T�zqn���xQ����&\q�� �U�A0>(�*�;���h�35�օ{��mtYZF��o��P�׍^Z��XE�Цg�g�똁���h�HF�ۙ>9ĪPNOl�x'C��ޕ8b�R�5,~yIfN �	�jN�n�FxD�,�JXSG<u1���L��`�dN�+Ȳ,��8�[,���xr�Y��I����+'�*�]������z�L��j/Y��~�U Ha�$�{MU-q�0[���VMZ��n
��<
��*2br����І΂����:�i�	$��^i�5��{�9w ����.��!O� q��' hCA�@��[�L��zgw!���jV�c���aۯ�R�/vw�D�\���7^���M�಻�;�xI��>�Y�v�0���T}�2D�Zb"�x&b�57��Pgg�J�m�E�Ƹ�9?,�N�5���j#�hd���yc��$;�'�L��dE��ۅ�����b8���#�\�)���Q�6��Ο~��=�ǹ&�4�0n�r�-���x�~��(``N^L�I���(s[�����n��빗\�M	"~�#,RDܗ�q^�FI���P �)42p&A��W���]OR��#V��ejv#�'��KOv"�2�.0��
�T@p�Q�6��s��d=�;lc�l�q;��JmR;�巠,u+s���g=>�%�Z�Z�r��G�&����#������~3x�#V�N�?v#�îoTvq�<��f��&N�<���4$�6BL����_H�ݨ�ǐ| ���I!���6h�+�9� O��<�iRT{�D0�H�C��8^���;O��-o�k# xjXz}��V�v��TG(B��',���ң�ƿu�����Wz�ќ;��%�J��XN4����['O��ɮk�ϗԨ_�YhE�1�:��|�Z��Q�^���ݭ\�'�i=�X���@x�}���t��Vh�XJiDy���}����1}�ʗ��>���-̳���&���>Z[�Qā@$��K#�%P�G�8�r�±��9!1��cd�J
�J�x|$-xI�X�Q���ЮM���.h)p|� ����	��Q��bg鋼���B
�0��/��k�yz�gN���ĥS�i�ߦ������ل�g^	������yEcM:�<[��Ύק:К����%�%x3u�M��e'���)�p8�ҿ� ^��H2<|y����4{5���C�7>���N�K���;�� Kߌ���J� ?�8:�@,i[�J�v*��vzUW8%3e����	(���՟����a�R�`��`��Q+��G�˾���:eO>�f����Ȑl�q�e������{M�K��_�����g~Y�3��g�E��[�8#�Q��sn�)M-2�
�����?��{�E]w�k�$��d6x�CrCf׵�*��g-��^�G��Aƻ�V��ɀ�z�0��� �Q'�Nӹ���y��u��u���|ID�( ���#��f����N�d�
3��DcI���3E,?$��W�u/�;'ɢ��e!�.Hб���C91�rQ��4x;6����O1�)����L��e��،��`'��N���*�F�4��p�3_�5-��Y@���a6�BKR�0�������1�(���$V.�ns� �z0l���Oۏ��8;�J�q���!�D�K��rCF
�&fH���X±�� �ԩ��AP
�3��Z�	��:�����<��=���ݻi9���������wj{0;	��0h��]�73Ήu��j?�J��a����p�����D�v�G	*�O� ����7e;�XUC�u�=ꐎ���TL8g�"�l��4���0WϤD���!`dR�'��
�����LuSn�=n�\�4�h��&�;[c}A�r��b�-k�f�tu�'V*�~}� +y���e�!����;H��5�IA-ǚ�չ��ZA=�����V_ ��p�3��"p��+rc��t�l�U}d#������]�"��g�k�]$Nm�һ��U�RtoƎ���L���������M^�J
��yɧ��<���t��U�g�&�!Z?�~VQZ�<�M�p:��K��ֽϟ�[rM��]��*,��轌�O@vs4 x������p�}��D�g?i*'G�����X˕��Q���eX����@=D�n��H�C��I��N��kƶ���EmBD�3�����Ƃ\���,�/vB��[!].{�W�a�=BB�J?�|��*�f�)�>�1D[����V��9��< ���!��`�c�6��֖�9!~y$�$H4)��T����-r�4)��� g)FҸ���LyrC�C�	2��	��ͣ�3zp�
^K��l��tf��oN�_P�l[u��#����=��^���jd�����Q~y��a���|M����|U{��xK{���D�J���C_04Al��M�H�RTl�_`G�l&�tc+��=�-����d��$�����O���
2�s���c���զB Ww}9�3��c� ZI���-(��lv�͓��G�.�bpz��z��8߅_�MĻ9�M���3��%��jj��s�X�ȕu���韯���R���?n0�-k����|��Z߁,{� Lm�Asq���h+<����:��So ��);}���Z�.;�t	�w�i��tկ�*.�C_����L�q�8����̜�_0�a�g$�_��/����b4x�^�؉x[n���L�d|;�(�֞��PLG^Q{^G��]P�˹ru,�O�ߞ1��V7?��P�o	�"�X�Iֲ�5��g��tW^'��WM�;���t�;�q�a��l��Ǧ3��D�1��ӽ���߀� 79$@�r�L�m&�:��j\8�HX扴�W;�z��AE>��v�xU;�J4�^����Ndmf�1�4)`��z'����>\����񴹘�����eH���/���V�T��K�M�B�P��G�8�ˁ�3^!�)Zy�^�Ԯ�j.c:a�)ļu�=��K,���<߭�N�>�2ޣ�jܶ���?)8��V�\fV����-��p��ePJ}�oy-�>���7}�X�ǽ�+Q����ܼ�K�@�|/��#� `��)��ЎM894{)���n��)5q����h	V����U*ug�G��cS����O����H eZY�����@�L��\�&�M4'𭕣:7J�mhK�u��^��f6��W��X�h+������kUX������R�\����<ʏ'32u��K�<򶼬�c�������:�Ef���g�5�1˶�B{���p�}����xz�V�?�Э�퀐�m�X�TAڢA�X��p>�^�":T�*Q�K�S_��G@��@��&t��Jm�������dK.,���;+X���)N��l�O4h	Mz���^�>,A<��$��5�ZCJ�a��G~1�V��8s������ʎ��|_���x��[�=f��]&�(��e]�9�{�L��i������72W�]�!�I!N�UZ�U�ɸՓmP�B*ԝɌ`�z6OiG��c���e@��饰���B�P���0��*{�$�~���Dt�[��\y�� �V�����s����*1넂�bQ�;������2�1io�+���1�A��g����Erq̊;oh�K��O;�������y|��ho���)節r/�v��O�{��y�%uP$F���`��D3o TI��X�ޙ^���%uX�Yڮb1��u`�"���H.��fh���Ҿ�5<ua8L �Ó�Z�c#\.���6���I�[�GI��WK?���.�qh�.@X��ϧ �m�?ڔϸ�4��BlHu6#�!QN޺(X�c^�&x��G����)����\�)�zu'��-�[(��R��y+�H�nf��t���&UNB�3�e
��`1BFjW1�N(����d�w�O�b]��]�^Ћ��q ���C99�O^�k���^/j;CfN��eK�=����[k�?������N"�k��0����(fjhd)��<���c��qmY�@61 ��#�%8��7�ZO%�N�ɗ_?��e�qS\[�2�5�b@��|���SP�0�E'K/d�U"V�[�ca������������!�o��CmF��8�y鲼Ű��aK��'o�����=����jp��b%���jgjf�D�~���ә2�O2�2 ��%D�BcEzK�T����q�Koi?=��G�e�?)\��(������V�ث)>��P�����)����+VO�:�m����xTp_#���H�@>y4�ٹ�\�x�RG{U	V�O��_X>�(�<�� �[_>�N���~��_����:L�:����W����
�.t�oJEτ�נ��l��W��L4��P��ZǎI�����jf^`����,�@)�e����.�~*�+Wp�O��6T��C�^_�� �������Tve�B.�1СX�*D��8������<h�Xvj�c�p0�?p�pXi@��#�\�d�a��PX�k�u͐������˫�t��SOp�q���ѝߨ�������+�����l�i�N����0��\�q��Xg�	�S(.����v����n���Lq������oZ��������[�j�ΪD�;U�u�[�c���IA�R]�]^����ڞ�,\h�mgU&�qp�9�t�Z��]�X~�9����������ܡ��F)Y�_ �th佃������R�BQ/n���q��~+�&��]w4-p:W����S(�3��%�ֽwL kӰ,8����2��;We
1��i�Eǁ%���U�"�p��'�TL�V�L�
�]l��>��8��0��Pg�%D����n��]h�ݮ{�0B�?��!B�'����z�/,?��q^d!�nOV ���z�� L�ǂRT�����7��[t���T�ܝ�[ٓիF�)�
��Z)��wR�b�L�v-���Z=%���}�"/��u&*'ҫ�C�a$�G�13�5�4=9�M�������g2�E��j�E�!�R&ҋq-�0dۄ �M�] %�>�R������b�@�lh�Q'J^`|<ͼ�����l��$���Y�rE��E5��|�0���W|h�Z���w�!�žo �󩊌�[p)�e|�fYyS4A��FrL�b0�� ��M��g*�^��'�{����v�kD�u�6�	���z����9�8o����7�@(}�x��E�O�#�Ir�
p����M��y�2���n�T��w���p�p��/�U~��D	�n��*��5{�p�e٪TCp�8=������F;v��:�c}�����d+�7|�*���I_|�\�:>����\�ʇw]i[�h�,U��vW��7��i�q/�''��w(��y��'�X�X�W�w#��/�&-��Xn��=kk)Z'M8��龶�NljW_�V��}vJ��`!��fy)�T7��֡�3y��\O��u:8���>[7[,��k_��M��߉`�]�-Dcu]��B��
?!�����#���:���e�K�~��R%^���k�P��BuM�x3�����O�5��2x�\�_�#*=�a]��H4b�W)�9k�S��:�O^��:�����,?�����ޤ�7F
zي���"
�r�k3�px�@}l�9b�4���r���c�@|1gYb��g0�̟��H�蟭�k�q��~�u<�qC���E5J������͍��E�/ز
�#!�:#�$�$��ȝ�އ?�"��-�`3xW�r�@���d:P���- �f�Xr�^�W��� �NRh�b��Ė����)��O��u#qT��l�6=Z����;�lb[��Q�<^ǒ�B(;��]>$ݭ�c4���	�m+r��仯��+�F��
�e��H���������Q�n�$c����;b��F�������Zq�ư-���	�a�P���$�+\Ƌ�tT��ц��b�\8-�v6tĥ�������As����� �>K*�6$y����č6���wT���U6�|��kq��ooKmh���
/B�۽��^/뵿$�G�dtP�jb�oqj�FM0�B8��_����I�v��b[DiA��|�K�'��n����	�]r���W��bb��>���5�˰&�5��w[�u��٣�@ @lK�H��JVϢ�+c� gF&vr^��km���@�E�"6�����8���j���e#���ߡN�����t|���_�PS/
ƤBn�����eN�_�~<�m ȭ���)^������T���BT���+�!N;ߙ���S��C����CM<d�%��x6��1_�=��ф��x�2�	
\���Z�1�Ϲ����e���}��q��9�W#�}����3~�jnG%)� �=&Kx5��� ^�Q�����m�_Zۊk���/��4���lC���O4ۢ��:](=j�x�)��vQ���p��*����C(�~��7�	�^2 Ւ��E��쑼�e-t�*��*$�H�s�g���XIX�ʇGѻ|����D`�8K�A�q`��lmdQ?�(�����%ͷ@'=��<x�{Q��c($�EV	�z�S���߻s�VU%+�@c	@�B�ؑ�����S���(�kd���D�*��|�f�sBdrD^���kW����������4�ҭJ�n5�Dk��]�{)��.ܔ��R��>A��
� �0o]��	 �	��.��%��j��2�Щ��Yaڎf���Qf�8�gBىP1��Z�+�.+��$o��:Ϧ�݌V�?���[�5M��'nn�Me4K��#G���
\I&'d(l�	P����tE��F؅,�6X��CoV�->pR��BwO��O�.N��u/U'�L%�)&Z������5Ñ�|�����}N��;_.�T�
��������Q%�]��l]� ۏ]�h=i+�ʒ�3أ続<L�\�,Ir�O�uVޟ)�d�� =2�q�)_Gj�r9c�yD��ߩ�����p����b��Iɂ���ᡀ��/]"�5�������U�kD軣r��f7�̮�K�(vu.��tԁ4�j�)- cS����fřr�"��ޥ��gC��|���O���qu�n� ґy�D�c;d�\1�R�D以��W��&��9���4�z@��}�f�#�"fȝ_P �fH��u��U����M�D��ӝ�}����y��A������{Ԇ��1.�Y�3��5IyG��������i��@U����ݰ�ԥr�hU}xj�D�����壵 �$uض�9~��c��r�I��[^��!m���=��z��/�٢��`�Ѭ������$�?	dZ:茯�G:|�7�� N��7�ƶ������="�@���r�F�AXsu��_��(2�2~Ϳ�,6�"�e���@���B��cR`�ТBO_�w�3�\\�1�2��I''�%���k_�H�q�����A�C��;i��'�Z��R��,L^Α�z=_s���h��-8C�PhK��6�_G��î��*i{�]w��t�n,���+ ��)��! o�ǫC�y������b�z�0m5�� 	�-�S�؝>�(E�]#Ks�b<)�-�2����`����:��G�����ҟ�`�.>̂�!�1�ս���%���eM�!�<8f��m�_�X����[��2n�8obj��ܲ��1�l�e��R��x�5dk�^�ઐ�������s�LD�r��Ud����ў Z��Πm�
��׈�Yv5t���۷����I/�Ȅ>�8m�"kG{���+lhVB��up!�P��7��W�b0[P�
���x�	g�=��_�rv/z��4{_}U+� �L��.ؖj��~�B���e�?��b�%㐃�u�W?�etoz��5r���r���%\u���=�\������BO�p5~\�wXйn�`¥*�tE��^cG+�{60��hb�� A�ՖB������H�(�:4�n�}�斵���rp��	܎�z��M�pk>�1D��ʃ��^Z��w3�٬x=Zw�㞼�,�u~�ͣ����+����2ʲ$j�l�o�|K��yWO��\���O���q8��o�fATս�S%S�{%0T�i8����g�ڒ�0}\�d���b����F�w�˿���ʤ������䱸څj��ۨy��%_��=g�9븋K��u��ݛ�o:n�\i�ܞsU��C���x��RD	&�M��������:�qUz���e�]z�g6�0@�c�߃-ф����^N.�9Xf�#����ǒ��TL��&?z�{t5�t����1���U�6�]��i135�s���E�!^� ���v���$+���#�u�WXow��s�:�&��ZW�8uĨC:g��|��/R��3Ь�U���F�_�fR�$âȕ$�P�c�I ��.�����~��5�I<K6�@)9o ��mX�k�e7��O5�/�)��V�\�M�ځ�Y����*���{a���ι|m�����#��gUL���#j���E%+}>wL�4)����&���ɶ������s& 	���52D
�~�M�X/�t����(_���"��4�f�l�6�b�Z����8q4G'
��f�&��D���	�Y+�����TvW�V^�f��!�$Q:v.�W���}�b���M���."@H��MZ3�s'�:XU��o.��`�����3�P%�"�s�|�qe��Ř<�����w�'c�3GC�qa|�^�Ŷ:�Z��s�C;*~oX�ȍ�O�En|�!�7�m#(yb��(��7Y �p4��7/ng]XC�	3��?z�F��o��ꄌ�>)� �ɣ��!����3_*�D9�A�dO�Բ�|Z� 3i�,���rf> ԟt�u`�(�+�
�;��RW��U�
,;r��~���=}?^#�� x,��_0�w����߭Q�V�A1e���4RQ@����U����[�:��cr��/S�#JE��#%K�i�h{ �J��?a����Sǅ��>�*��+;t��p�>/���gP0�D�@f��qKf�J2����e�����E��ՖB���`FX�� {�Ԗ/2�tq��)�\���f�][�l�Q�i���+�44P������v"�IN��z��r����@�^}��m08�}�A�>(�zW��Ɖ}F'�`)�*ii}:���)�
�5F]��|�Tև�ر��r��ޫ�����l��j��+�*��8���� 5|z\���vʞ�)J��טY"�(1�5.6�5#���>H�G�O�����}��F���-�������њ�#�ٹW��W����eiJ��;��:���#�zt����d��]N2us���a\90�@�)�F��"��\��/�|��++!3�B����C�Z�����{�����;��'҈���ȼ���3����Y9m�m�k $1!Lܕ�'U�-��՛+���,i\�gx��5h����L�b������	�� a�Z�#ՠ��'g�c��E��W�w����J�]>����L��<�>01�Ej��by�&���h7��?e��\�z�ܱ٭�x��Ӱt��i�J�w_�w�:��E�e�s7x5����eC�-�n4�a���>��㟮W��g0F���[���i��'���m����)Wv�V訝�Ɓ/�6�WO�ds��}�t��<�,�SB�xK�C<e�7��"���E*�C�����^�o��nCU�+*�I�?u󙥯=���A
��Ο�JO� � C���_Ǔ�똠��fM����Kb�En[N�
��LՊ�\Ky�P��J�P
F��Q�1�J62+�I�/P1 R�n�O�2� s _� ˟F	�Lr�%��K�)�WG�8�8��G&˖��q��Ǣ���:�^;u!�/��ێ">&O�Kݟu��[��sU ��70�w`�t)]6����y�ig��n{
���R��\ƨc*�٭L�)�1*�p��9��1FA�1�����	�-B����Qx!6�����Qڇ]rL����"�����V������IW:7/��#��&�,���"���"�YՖDQr�=I������Cd�l�� /P�'C�bC[����4�1X�9;Д��w����c�9�pt#��� ���4�G�#��J��	�p)G <H��N
�C�-3ڔ����q�M	�d����o�?B�#w�J>l�x�d+�0�D h�Vvب���@Ʋ8������ɳ�nk��~V��.�ވ��>�nد<t�v�.$`�7	��d��x��%��RQ�������S����A QU�$ )�A�X#�>$5�B��
�9N?yQX��VBWuUf��~(;+��C��������'ld܆��y�`��gLʩƍ�o�����?am#��3��k��,���DQE�M�n�֗� czz��8DX���AY�X�k{䪡)��f9�)����/�Dg�rZh�}H�C=$JC��n��^=�>ϫ�T��DgDP_����r�
��4��٩�tҞ[�G|A�0�Z�ߨU�jb���þm(��B+{��v��b��� �6�ܛ�l4��º�IS٨~	�7�N������I�m�j�H�R_�8d�38H$��B�f�VbV��[&���5�l�Jj�q2�9�!��{��ʭh��q��}���N�9�&v޹�V���-to��}�n�"U��$d��oP�ϻA|�<�"�4�}{:��į�:��~41��Ӷ�E_�*aF�<u{O�`�2Z��~w&������n����Q�D�>w�%Б����l��/CHn��->��LT��cW�l��{��d'��q������q���ZdVp��F�9i�i��t�XIg��Ȥ�����j�<�Y��<�#0�D�!�Bo�(��K�Q���~ח��Be�l�1���O��pVH��0�5%��>� c�F��]��2��N �;�!1�	���@�:�V��4����GZ��^o��Q���� �Ԟ��rō��E'�u��Ň&�$m~Wcm��q��M$�2�c&����s,����x����Z5���*�H�c���V~�m{���Lz�b�n����[N�ݽ�k<�l3�tT�  @�R��5����!��}�M�A�~&�vρ3DLtJyc��j�d��I�,*�]a�)�K�t��}3�W��[$�^�Y�r2˶�S`����xF�|����®��QO�K����O|�{�MUO�h�t�l &��h#��]v&�J�+ˬ>Ы�L�
{���ά8�;���*Y��D�_Y�;�%Z�����s�X�9�P�u�5���P����\�,x=p�������<� ����2]�7�3���a��KY"�Q
t��X��B��^�j>��at�Mrb�wA#�� �g��o�3d���p�lQ�9�35_�W4�)��c���Zlф�9=w�ާ�)���l��Df������6�s�Ǚ v��)Nӫ,��G�W ���
@U�'�j��fz��������	�^���W�.A.b���a��5:!<�s��im�	��B"�-к��`�~n[j�c�j����u�T�4�$�������D�,r-Q�8�W�1�A�y�vtUd�Ȅ��X�El�m�e��������S� ��^�u ���r;�?����r�����O	b\��R��������J©�7X(�z��Z��d�i����M��Z
����(Q���� ���$;4�o$���}�n��V|�,VuX��R����|������h8�KS�(�<��)?�38}���<_��XY�|k¬�6��a����cr⢦X#��>@�/��hQ���\�~eUxB�`�a���Sp�ɻ�GnD[k*�n`����ٺ��=d˔��ݗM���K���˛���[R ��q9^��)��y�8���.��Fn�!�vL'{���֊���pýCh��24b�3�������߄_ڶrFIBƂq�`H�ɠB���h'R��x�P����;��� @hb��-Z�\�R æF�:�t�
_x�Fvc��F��X{�:)���	��FӯT L�_O��dT�F1�E���ok�I��#t�X����ڿ�(�9&�2��k4=��I�I5T���F��Zw��V�9YM+����)3�^~�L���d��_7�5�Fb���w��C����<���?�˖��$� i��l��co�ʘS��Mi΀Ch��K$�n�G�KF��i�ˇ�¥�|�'��������nG/��I��X���t��kC�<h&��v��j��|���0�0�re%�����c2hTl'���߆�/Uã�
|���X�P����tzP]��B��ĳ!!e0mb��>�7�3?x9�VS���'����6>�K�MxӤ��Vj��Ͱ��a2v����1�!!C!�`���g��W�j����Ϟ�<h��0�;�cN�Q��g�>�1����s�nA���V��E�zd��ÃF��B@�3;N��Pb�!�$3�^��ifs��Z�&����)|�A������GYϨU��Lc�%9K��Ɓ�'~��M����8%�
������.�ܺ�Gb�Kw��8�W�#*<N�`����Q0�1�QVk����Q��x��OÈc?�/�߈w�:[���Ҷ�Vs�:������0j�)���^��O��+���Ҁ(�K�s���tU/Fvg�K��3-vdxMvR6Ȉ7^IYUʛ@C#?	�{�F���n�V}�CL�p)]�hc��YA�z��(��M�_.}�\�K��\�q�{J�(p��B���]k���v�ߤ����r"ɔ����\.z�y��a���wU͹f&�e���]��~F��1���Ȳ�`�y�Y�1x�zJ�`r ���.\��[���<Pv�pK� �7��mYeE�X}��J­
��{����
{��
��hx9 ��kU��  ��n j�{p\5�Y��*?�v<�����Fx4���f�h�����ұ��쏍��}�D?��{��&b98�]�C���!SM���.n�R��B����%B��C�moD;}ѐ}1Ř���*��+p{I7���u��S��$A���&P���X�Do{ik��tV��j�����)�3���Λg�pݑ�z'�4�̊��3^�DL��������]}���k{�e����9������2��i�WK�V�_%�Y��;�ލ|����E�P���vO�F��I\��6I��������������y�6�#�W%h[��:=.����- �=��B����d�/mI��Ԁ������`�V�J�
�o����4��>��cf�%+d6�T���v��F6pE���H���|��bf�	�R+xv����l-�Q�p^R�j(�Z*�M�1׍���m�����7�0C�2%FK�%�&�7���yD�́Zj�Y�,���n�uP9zmvQ�'N��+�@T�?DN�ri���*ș+�L�Ża�ƿ�]bL��saTx�#�ɇ2Y!��)��wC`��\��#�&��)���/�#W�(`ͫz���O�X>�����$��!��W�ʗ�_��,�ޘR]m�,�~�jK;���9�\�A�?tp* Ҕ4��t�1��h@�qU
}�

h����:-��u��Q�|�ؗ V���s�^�x�
m���ən���nXڠ��L��2����Q�;��������n�+�����9�#j���À��1|�I6�R�z]R>�!��
�i�YLSg��H�
�X%o��j��ǀ��Ȑe�Y��3+�#��L$j���,�'����\��#��EM��@D܏xY��[.��j������3��ʹL��-'0f �>��c�� o*��Yr²U�㉍�!�,lcBD����]<(�8��㋍Է��,аP��S��
�iL��\cV�|���b��<_E��n������څ�˅Q���~�,��ނ/!�UʸO�L6lU��D|CysQ69w��}�F��0gkp,�{�!��c���Ƚ.!�C�e�y�g"uO<�k�:<�ߘٕ���ϘH>x4��*aK�1�H�wh;;�O"��O<���s�/^R�и�v�m�7�fv�i�E�i��D�����8\�&��yu����Z����8Ů�K�����������)����H���!nY1�{D�A�O<��S4�����V܇�I\��ӛ�$��Omx"��c�����՚�-X&K���Ol�64!�7�Qa�X�j��>Bŵxr�vU��3lYD}���q����a�J�{�?_^�����‡��M�㊨�;��?>�#�(�P������]#�z	��`��ze�@ϳ�����\ڟ��\ꞃ�%�e4�����a�T��Bl��o>?�ź>#� M�/*���u�~�c�8�}g�'tVy_��S��ù2dBR���������;�'�Z9���N&�䤹��y�nt|�~o����>�'
��*BD�"�2o��,�#�)l��)����(��981�����d��Z�J1�Љ�L�EJ���q.Q���v+yL��;��:���<_y`�h��4�`A�)E�UD!�}���`H7���!����s��aʃ��%�>�z��Y�����N�ꆕf���=�d3y� o�{�Y�6�$݋��|m����/e�9�����7j���IkaIU��~`��Ig�M,Y�s�E�7a��n?���?���ám�A�q:o�����l�^lv4�LA�\ �0{=�|��a�w� ΂8��=���i#{�ΖT����c�ʜ��.]|Ț���q(�!��W:��G�i�A�!�a�ۿ���t��έ]2�R�m3V�ǌþ4�Pw��Ή��Qd
�+G${R�#L����El&G����ʦR`�;jȇG�S��R�	�)�Ry�+9��fu�Y]�sBc�,1��pO;_z����/TZHM1z�Y��ɵp��"�� ��[{.�/��X��˼��(�W�؂�?l�k#3Qc����0�]�u��=Ϭ� g��.�E0Ѱ�~rP�G�Y�����,б ߂�r2��6&���GS|�z.9'��Q$��_���&v#Y�dת&w�<��\�Sل-��w�A�J�所-)���I�0��_b�"�D$Sz��ޥ��NOOڠ�M#��Z������f�ޘ�N��vJ��t�c�T,g��_(6�轡z���fU/ƮO�8��
�B`�� ���!ѳMjW �����4x�]�y�5hm/
���Ķ�B2�+��+&��W?B'�i�a��<9{#��n;��֊h?��L����->�k3��E]C�a=F��)�LF��+iޟ�xF�V���^��y���wd��$F�:�C��l]����:���tg.�F�S���x%7jZ��넝_;���y�u��1��=�������ס�dm�k��\�jN�Ц�%n����	��އv��~V�
9w+��&�O+a�PQ����u=����!��p��������?"���I*��}{�V,#�Z�3=_�p+ש�T({��G��,1�����M�j����.a��������}݁�!O�_�y6�����NY�g������u���{w,��H�nW�X���IX{�_�MSD�qAk(�����U{��:�=�ʜF6���#��}?o�<��`�rL4ȱ�C`��t=K�O�^�����ҡ+��1w��$�_�C��!�սs�d��!��0�9����a���"6'��/>_I+C]�Is������1�0��fC�[NpD���j��X�!u6�6Ps�,F���R1����v��F�o]&x���b��j"j
��0��_AV5t�٢q�yk�������������p�`�7�!�M
e��+;��+��~�|��+O� �}�
�i�Ĝ���	e��=&~���A#�����B9G7�m�pNj�;���=��l����.�g����s�/y�}��KDoZ��J�*�d"�ULУ��9���1����e�QL1T�XH��0���q�Y|V��0�r}���%sU@�9��DYD��Bu���)0��t��������g�9|!ѫ��K�ԛM�>q��������ߺ�����R`{���61�h��	a�p1u ����^�s��n�Nu =������g���>�6ν�=�x;��B�>%���C ��0Ab��RؾT�
~����� �M�P ����1�{��!o]�k�J-᳹�ef�I�Ilk['KC8�]|�>Ʀ���ޯ*� �$�d���,��p�JܦŃq�w�'�A��
���٩1�;��������]4�x�9(Nh�-�V��)l�BE�3�����_�P=��V.���v��a����
3���44�&�%�g���U�[:UF&;⏜�v����R�@�A=��g⻖���[!+̢M�_y�������Υ���r�ٌ�rl�;V����!��V쓷�L���|�$����&�ҰpY@Y-��x��w)Wޘ�޺�@<���NO�-uZ��j��G�����Z:iz���Ë��	 �Vq��	˄�Uh�^0��šW�3� ���z�T��%��=���uTe�B���m\(�q��3�L�	&k����|� @��H@�Bb��29�����n��p�VT�1R��Z;�*�lT��Rkz*�	?g{#9����&/�f΀(b5�c~���c�K��*+Sz��L\�'����?�U����Ph��ur�{'��5}U��>�����VM4�"ņwxYk��'�Hzk7d]%8�gpJ/�>�2�o��,�Ճ�EQ�F�ޕw�,ec��v������ǵ�wi�ژ� QU���>�"7�h')�Ⱑ�Q�9��%o$.���`m�U~hv˵0^އҫ�^�2�)7��m�ZO1��j�Kɜ��(���ܢ�4�h�:8H�L��v�~�F%)L;_�-"�\6����I:���=ʺ 0_N�4�M����%]@I F��qК8�^ȄM�^�ϣTu}H��A.�4-�����5���Kϭ��7%�0/�7,G=�L��B����Zt�x���f%a��*�(�x��DH�5�]ҽ�ٴ��+	����V@���Rm�����r7�DZ 7�,K�5п����X]�2�NjC��ȩI_�|,τ��eA�t�`��S��Hz�Sß�k%��$CBp|Ĳ�N�H�X�{���؇�K�2Б1ȯ�M�(����;|-Np4i���ceE��b��\+hM�%_Vƚ_iB���j���6fK<n���6g�^� ���[QԒ��C\<�?Z�����_�PT[ne�'�#]�X��	��9Պ_�)�.�ϟ��
?��z��B���s�O�>
�a�E��2ݼ0�p��.3y�q���r=�^���%�ޟ���s|�&q�R^�I�ј$l��zزQ�h�&����{��j����E�^	s�YFoE�cn�S�kv�/�9�*q@��_�c�;��*��zZ6�!�}�4,?�:�\&g��K��@��c-��*�D/���q�½e��|FK+X:�����Y�K��QeT�/:8�،v�>�{C{6X�M�n�����;�_:�M��0BU�t���V�n��@YqG�姱����GluNW�,ޙ�ou�L]�t����B�v����|�\���Yݹ�jr�_(o�f�I�T<��/C��,ZWa��8������	����t�Ũ]a�W�!��bV=� )(Wf51h5�Y"Wu�����(�`"V |`;�%^V�0a���}Q)����lɑ���	S��8�h�N��y��5:�e	4��ot JÔ>'tLF���?�p9��ERl�di�F���'	�<��/DU������^QM�9�_����l�B�Ři�*�4�M��zSa�cs{�C�K�r����1���?u����U��!����κ	Ԡ�Q���T_��͓3 �ׯ{��.��b����"9�6z�����7;|ڢ3���"D�E��7�O�kk(��s�4�*6���;~�#�\@�p���vl�:�:*���Hq�5�����aWzd����3ɟ���Y�xX��o���@Je0�C쨿���6�nD*s���5�G�a�A�帛�磢��I��mw��5>�x��Ee���Ьy���BWVBo�gN�U@q�Yh��Q����=-ڹ�@����̬M~�"�`�u#��
>X��R�&�C�]�%��ӄ`=�,&��FSevL�q?�Y�b��&tGiD���?o�e�5���u�i^��S�5J�ٱQ���7B8Xsgiwu��������v�H�68�Uw>b��ѿВQ��,��%��������������|dN��V��G����٭\��L`��0c�x8R�?&�2F^��˥[�r	;ӌ�}g�����/B�1�v#ҏ�=��A
��&z����#�ݜ$�15Eql ��s���ёTNt.L2�^w̒�g&���k4����O�Ϻ���aa����#&S��M��G�#���箟f��p�o�%�7}:L�H��%�ڃ�kI�Q=��k��+q���Zn��f	V��!���ֺ�㷐vVpY$��%�8ԩ]n�ɻ[L�˫?�� m�'�d:*����؛��p��"D��|<��?��_`��1F�������?��W���}�Q�̳i[FX�����C��.����N9��E]�;����h�VQv*D�ؘd�V�B�[�&v����|=��o�Q)I���+F��zN�gxR����uvJ���W5r�Jj��S�%w��s�3, +��u���>���}EHw5�W�:s����7��<���n�&�=�Ԅ��*��\�#��T�T�͓f�N�g.�у89�FJ �Vڄ�5?l�ٯ�a4�
��.�u�S�0u��FJ��-�M��M2G�[WA���5}��F��#�4�L�i�ҭ���h_��GX��W&k������C:��}�:��X4��ELV��*�_Y�:�je^*�z�p�uխ�gbXXPI6o��o�_��ܒs�Z_I�_f�CSc,
�����K;�֗��56ӿ4�D��ZV.�b1��MizI�nL!�]�J��qQ{Kc0��ʓ���ї��
�G�#��;��)X�]Eh�r�i=�Y�n��D��/�UN���Vԡ�V`W�z?ǍK�C�G��W��t���Ǜ��s�UB�rq�B��Wa�A���Sdp�����-K��7���4�~� �ᒕ�[�y���V�!���"11g�����F@	��1nq��f��(W#�G/����J��l���8W!;л*O�~̕+�����s�p�_����:Ⱦ׽Gq��dCKo�'N�k^�� 
&q�@�+�ҷ���Ġv
�T�3�Ip�������pk\Uf࿀��q�"�4�듵�k�,��A�H���,�7�,�B�v~�|�U�r9v0 ���`�1l%k��LަjS����޲��GI9�ȇ��8~9�pcb���2�muɩOP�ɡ�Щ__�f�g�PD��n���7-����Ԯ2E�t��z}�m�d����4���K�O���*uٚ�,�T��a�rN��	dZ�	ęXL�P��:x����&s�8�iܙR� v@��K��d��t��y�v�
�d��&r�9"RIb���-<4m��G��h�xnFh�����~rX�ry��
z�h�/I��$(GKoK����<S�7A��m���BRS�b��0�k������� R�-ЂZ�8|��.�Zh��Qs��`8�-��ݲ�S���>�'n���S�b�8]��r`�"����Z����+bk^[=7�NH��"b=���0Ok�n���W,��Qj
�]�5^Y�8l��e��{ �ܰ|�����		w�%��ՄD4��^���P]��$k��d1?n;��;,�1�z<л�@�`����r��\��M�r�Ŝ��;���=�6�i�>\e������͊�� qqp��m,	��Y~�'2X���S)m��KqU.'���]�>�c(>H�E �ۊ������@�d�遁K�Ǜw"�qH�)(w�G1����n_�ʉ���R֫��8Jگ{���"��W�(�r�lE�z0��rkG�%�5#�T�<
㓗d�����=���b^y���zoX%��	�e�fDп��v=���o��8�-j��+�������"�7�{�ƬT�=$��Sܔ���@�(�ҩ�:^���L@0�IΔ�?L�ϩÇ�{8����dF��#�A�6�
U!�	�X���?�.�)v��.	e�q�ϝ�Z;���˛SG���u��kL�T�c`�wZ��Q��d�%�;~b.�d4?�0�~!T��'�����n�R����.-�,�|"�c�`A۱M�+&����c����ϧq#�ʜڌ$�\>��kz.�듮������<�?E��0���"8>�1k�ʴ����T(�Q��y��q�7�͕Ixd!�ez\/\5T��"RoO-�p��RYI�x2 �d�����@���X'Nuv�#d�	#1.&���������{؝B�������Uc`���͝Ǫ��߷��G� .�T��w���e;� L�.x�'���o�`��҅r�o��S]b��$�R<+:w/}T��J�7z�9)�O'n�����	'A�N�W1��;��D����0!����S8
��M�W�c�K�o����K;���9Ҳ��Ǌoe�i�	�*s�aN�tB�Bo���^	0@�m�+{[�_6g11I��=���l�|�$�u=>��M@�ڐ<IT�]�F?��ٌ�$	�	3@�z�������  >��:�L��+W�"�ѳ@Yѹ�d|�A"�Rs�DT�ˆA��k���&nY�=�����,�����������	�R�цK��5�� A˸ّxO�/m�rؼU��CgBZ����k6_����&l�kT�0�j+`��1��)�F�brZy�Y"6U�����
�����h��"K�jV��ۦN(�c�e�s�r�y[�=�ʜK����L�����#�����pK8A>�D�#�ʛ`��Ԓ A�2OOgq��!' Y����Tk(���\��y^�qT;���O�gN��{3�(KF�"��|~���?~��{3�9�m�{�5[������.�c05&�^��V������Sy(����ū��t7��=p:q�+U-���6o�_�z)$�:�>6Rk���Y�R��)���*�.ے+R��|F[�i��Wwrb ߔ8{�*2�B���Nܴ�!��{e�|xO�3�9OĲROͣ��@�����q�@>~ꆜ�����9[��kR�˽�F�*�o�¨��x�0Via��xݰ �ܥ���e�7��|Nҩ�"�8�C�/��J�PJj��y/S��x���+2�z��-�� ��'O��5v˥.��@-Xi���t��ګ?�����E=o�A5����,fQp�d�O�"D��q��U��[����5~��/��J���MG��._Z.���I9�����|�h< 45�%�1���E�3��!��1L�`wb�,*:MK$���Ad٨g��H��5l����������k�eضl:38Z����R�n�^s�̚`��IdK�#1��- ��e�w�|4]|��[b�t@ʑB�$;c
w��Zt-��/�om�k����
0:m��=5?���8�ޓ��&�����^�~5���-������(�	o-FdE����m#9̄��8�꼡EM)���A��HQj����@���HSx�\�I�ke�?�RK'w+� SQb㼏��b��7��d@/���k�{+@:/Z�9�Yt�S6�l�� ���oQ�K�I�;zW�5hS�7�<��LY�~4)h��0t��~=	0eW�13�j���������0?��];���ZMw��r����\����,���`i+�G�u�x�6�l֘��bX9PDx]r�������K����k�syd�6�5�Fy�/1�w�[��s�(zٽ�Ӟ��PZh%����U)��{������'�c�ע���OP�R�D���Q?>�'ed��-��w3���ߗ�j��}˅�S;hU���\��Ú�6z�����������g�qf�yXw�A���\�-.Y�,7(u��l&�4�zi�y|5��j�H��.O,���3)_�pb/|��$��p��RY<	~%�dTK0 (��X��%E%b3��0!^Z+�^�NbWc�����)�~P���`e�?r������b�y9�|���MC���.fO`-�V���Fe�X�{��1� 6X�
�
�)���.��|gMD�P1�n򜃶�UU`������g�ago��Q��B�~R>䄺��P5+�(�pӿ�����BEC ��Y�k�.�T}��.�M���?I���X�i�W�i�v(j-��X���9�z�`&a��/	纎�5�TX;k\��	QT��D��x�'MA�����C\��ߥ��[7FU���S���+�+<Wg��[}����I���HQ��K��[�S%���2���9���gyr�1L#����-��N4O�;tWc�^�/CX^h��,)��X���J�0��^f�.�ۇXR6��2E�_���SO~����$��ϐ8��{շ�x�j�����Ęh̵8!R�~���n�_o�K_Pc�m��0u4Y7�(t�}��o�bEr��p��?�Uߡ}~{ ���)��<������~�'S�(q��o+�4x�������6���� ��ξ��T<��/�وN
4�X�q!;<J,����ظg7@N�'+���-�r@n�K�^� ~]�<��<�U�n��������삠|�rqK�!9�n�i�˵��W����L~ny7�=ԭ�;����`\��?)���h���������{�%@��ϬMe*���+�5}tf�מ~PZc^G�	4��- A!eꩇ=j�����B=A��<\co�*�p�S��8���g 0G���j��q����'`��lfS�NH;`�=P*o,-��0\�U*pЪд�iU�t���)a����ӑQ�*�G�^S�,
)��jw?�4m�H:(Z6���\��,�P8汳�EG�T��d�$��am�CYe{���؈ـ[g�]˓h�ػ��F�>ޒ�=~�ۍ/�
�O�0����jb��z�9��R�"��(Es�jv�qH��O*�<���h/� Ԋ�ҡ2��u �QL�5>> ��$˷B�-�v��{q�[���f&������h
%+��4�7f�DU�m%"s�w��)��8,)g�Kc�=Ȃ���>���iP��8�.?��Ħ��HkZ�>�%��v���r�ߺ�;^@|t��W�W �K���ٲ-
�-�S*<��fl1��c�:�#�9$!Q�b�� 3����5��߈�_���������L]��l�h���fDo��G�<i{� lCwV�������%SW�������k���؎��tSc�E(�g�%חwŐ�p�� �nW�����"� �̏}l��7^�=�c�%������Oȝqm�d�T@f�|)72�RQ�1K���	����}vt��	Z���8Gpq�X�Cyd�t��AH�vBUT���};�ԗ�ؤFc!�\[�ID��3�e�����R)3玭�s�=rU1G���$��9|[���ky��#�3��-7��a����M4�F��6��7)q�?/��:i��\!g�1GP�uµ��=��;N�T��H<�(���=�����3Ė/y���~�GJ��� �$��|Oς�=�ӞZ��K��C�!^�����Jd`��xYat^���w7��v��y+�,iвWX�3�}R����6P��?sΰ3����\O��
"4�3AX��&��1\9�?Z�sS9b��`Q��{�<�t��s�ٍ́��i��A�[�78}t1?��x�:p�#�V�zJ�jv���7�*��^*H0�6NHj;}����+�)�	x��(���(��#�`�Q2Rk�>��,NG�(��>ܸ�N:ē������2�e%`?Y�:7+�߉^\AB���j*r;D�d��/_��[Ͼ��C<{��zeEÓ��c<1;7�����(o�����h���'!����&�X\p��D�AK���D��}ت{ϡ��Ɔ�g��0%h.�Mx���9ڝ��@2Bb2`_�<�E��è؉�5�[��Hܤ�.��Q�L���8� W��'u��K/�7��o����t���e���8�>�7�?k�P=*8e>��(M��'/q�DR7�Ģ�`m#�V��a〈��ZJb/�[�k�p�ç��$y󓝬Y��;o�)��5���C��lC(������5���]X����
��������ʱz|��V��m��&����a�[��e	��e���m�^ C	Z�z�&p�?�J#!7�K:y���%���Q�����P�8̉$���$n��u(�����U���T���:\��n�\h1%8P7G������<Kj"4h4��csn.���F�sY���4��fuZ�_k��/*zE��!�^f��򔿚5�#�0"���`s��Ҝ�[�Լd�
\A��"�� lB�C_l�i��⡭�I%Z,��Y{�Fy�G�H�4p����5x�g���G��xA4"������/�櫛>�O
&1��;۪h���Z'f���k}Œ���lzr[�-�G�`�!�2�o��
�����_A1G�+�HZ���)w��u�R��H��cSd���!�N�*��սy-��%j5/MKRC����bwiT�~(���?��b|a����fy��ٹʰ��$�jj.���j��ê��5�G�W����c�#�fc@�h�[d�(���E��g3=E���;r/m�]:�G\�AM7WO,a�uT�M&d1���u���?��qm�0jU��]�a�"���.��e�CܽK<��4d��	�
�����{�����U��V{(�s3�R[�HS��o)�G
�.�������k��J������r=.�Y�ݾ��F=��J.�d+S	�FG�:q�j���ʷ�ޠ�������P�˗7u]JOՙ�پzN  ����UY��]�|��nο�dMu�����v`��A�y�˳f��(dy�n�>d�R�ʮ�P-�il��S�R~ʐ�3cI�CjB�20;�6:��B^�:rL��7��L��4~Yв5ׄ�i�D~�[���Ho�qsܘ���2�j��*5u����&Ja�̿�T��n��}{' ��K6ʞ��1EP ���7�3�2�܃�Bl�OE}�8�H�yVb�a�苝�4��I`��D���͑C�A@,�����qR9�n-Z�H`�7�&���q9��	�y?J�e�a��c�a}���C��Dry`n�1��[Ŝ�-�d9I�J�ܡo������V��N�St�2�N�!�qc|�}ӕ�bA�ޒe�5I�{m�ﱦҿ�rS�A&Z~��U���a��Oet���.({�D!9f.����{/����!�h*��8X����6��@{���\���:Yh/]����xfů!�{����O�&'Ny�)���l����htq��*�C��e0�F�^��>	�.�9�Aά��
yj(�)`a�En-`�X���6�&(^Twv��Dgұ���@2�4!�m �%����'�4%��њDOkx���go2�ѣ�J���ϏM��.�v�Sֿ�9*ᴇ�^���߫-$���>39��v��}���dro���e���ɤ�`�Mi��b��ErZHr��W��m��f4�s��<y���[)f)�1�c�m%�E�!�=�w-����i�)��;�l?TY�
DH����0c8��J ���;`���;�p��24O��v,5�sA���d�Y��wzJ�;��f���G-����õ�a��#�!]C=�+�BN��R�& B���Q 6����n*�������0W9���]i�C��y�0_!\�h�8M��87����{P�e�4*�]��܍ _�� �[e[����"�րlh��Qr�`U9�J���j���R;.��oUZ���M�6��zɃ�Ů(�P��
�l�Q*:L��8��'�5�0^m9���ϵo
#��:�fa��|U�'��X����L�^��e("�V��>�Z�0���:` �AP�/��X̟w����W};
p`��$�|�09��Nł�-k+D���v���ÓM%����Ӑ��^�7"�-t�lt��,���ݏ)3w��)H��O@,	+`���ކ@Mp+��
�ZJ�91x��{;p�����<�|��C����sn �{���i����ꋈ4K��F9{3�%� �;��edʣ��֡���+�� �Ρ�X ���	b�E�k��r�w�&�Z�q������������pd��t�mH}sX
�7��xU����\�k�;�C��|ɶ�7
Cx'�;�O+����o����c<Bg��WӨS82wǏ��JO1�bw�~g*­ �@�0tq2��+.Eǝ	�ɌOm�����#�gL��F�3�kF�zj����a���,�bM���4��+�D�����y�f�/���C/E�
n{&;����D'ፃ�s�

M�r�s�w�?�����.�U���z|��9�F&�N�c�59�5�M���_^;�T�k_Sj`��0��
�qD�&��N��c����� �#��ہF�eJH�z��=�J��
�8�8(�4��I�\� ���(v��hra'of�4ԈVz�$�����)�,z=W,`o_�[F4$U|�wC���WGA7Cv��l56p��bʛpE��6?\ᑏ���y)lbw/)GI�{�gt4N�XҌ��n�����B.����黤o��R��T~�І�#PoG���tY8W�HO�������a���ď��\���=�J�=;�$�Bj��M�If����{��.�`H��zƜ����D�}D�S�[�p��ۢ=���z��V�^�d.b�Fݨ��yZ:���,I���QPӪ�+�.tFy�ڣd���c~Ĥ��zE��̰p���k��ZBF'�N&&�GF7��Ȋ����~��nu�jy�v��̻�~U}�u��W4�h��䱗��GĠ����-���'��΂��ɗ��һ='j}ڒ9��AӠ��H8�<}Wd��B dѺh�"�IlK��ڨU�p��%iĘJZhp�f�C"&�PR��ݾK�ĥ�n������50�&run�C�H@�2�t(�����M�[k@�-��/��8~�=����Y<:�r�&W�w��L��h���b0�}%ޤ��֥n�����qҢ�����Z�^�i�1�(���5�n�ǆ��C��JJ_�m������F�7����:�LD_�ܡ�4x�Cc��9���;�����4��ק�ߧF&m#jUM�ރ�t Mԗnf��>�W���s��cw$.����q�m�x�u7���<|uasv���P$�Y�b�;��ʝOkI��C<#�E��D-���D�q�ڻO�N`��4g�ۅ�8a_����ċ�`^�Ԟ�?#6N�yjp`��s-f
�Us�U�]�Bi����4����߼V���ox��j�׮׭L�u��H-��때J�� 44L�bo7>��-��h��J2���4̏gv���k�O�زSD#��� ����,ߪD�DyI�
��I��	!��l�x�Bҝ0.�����HS�[��}X�i�g�UD��>��D[In��L��Q�E �s���O�5���:�]&?�\��|v�����=Pqc���j���! !���D�\���tcU�f�_:�-ψV��������e���/�ݣd(�@_o�wr�^?������-5��1a��`	�qwQ���0Q�h�|��#���W��>��
�y򁋟A�_�	Q�$-8��d^s��X��J�8����ߤ�ZR�UI��s�D/��v�����Ŵ"/"�V2���ƕ��U[#2�\�5�6`b�|e5�(���b/vf"��]Y��\�� ��P���6��
����Kfr�8
�8��u���hb$6{̥������%a�LyDx<2Zb��g����d@(����=䅳Q2e9_���e�ɹ5�����թ�b��jq�
��7�GP��`!��Nߚ"���������(j�ɳ�e��tp�/���a �2�8g�f<�w��X��I��������\��8�(�Hљ�J?L��i�.:jP��Լ���.���}�4���OA��8^[.�S�A?��D��).\��Zf�{x����2�^k�|z\{T����%�Fȿ�9y�7�neL}��n��OnDx��)���V]̈{p��Nd_ߪ`-�ǟ1�����puZ�[�����7p�U�6T�B��*t���?��Yf����);�,��'�4�F(Rƅ-�5��'�����{W:�'� ��tWK+G$Sm��|�̯��Ǘ��O����	�����(��~��k�Uȳ�qE�K�y����B�������o�������z@��z�-Q����2'�ԻZ����ltթ�w��ie �
1�j��!:���2F�7��ˡ�A$x9�۶�Un4N�<���G>j���&�<�+l����0�X���*l��X�c��jRL��T˙'t����\�/��)nσ����VzY�}®�^�5P�E��.xY�׎��yh0'��vz�OM��HJɫ�V�B�(րq����i{��PL��y%�k�:#K�M��-?����ڶ�< ޹�>h�l� LHɖ���VD]b��@[2w��\>�b���ס�����^�#*��#[��6�J�r���L.p�xy�v��c7c������XQr�}Ղ�E;�co�YK���h��V�/�{C�#�k�N�� e8Ԟro�u��R�i�,��~E3��>�&I�	MG�Ō�Q�1?ŇF�����7?p:w�H���{
9ĄV�ڵ�[�g�8��,;8��=��k�=
�D���h�K�E�RB��y}�*<S�$}���&���	�=��&߯�?�v�Ț�����Pz�P��������?�G�z��z�@��Ш7�</?������	��2�n8=�n�K���q�ꅸDY:^�����#Lߏ�њ�'��W�+���$9g�Y���C���C2�1�{�
r9T�%��;��X�z�a����[D��ˢ�:��;{ �tm/:n���z��]f�������fg�ҁ4�#��R)^D�:��t��> 4Y������ϰ���x���Ծ��2tK�FDD���E�w=_⌏�m� �֦�?��8�����W��
�x,jk@�22T�E2�7K��osSD뵬֕�@i�Eo��\�D������!���PrNC��N�:��j��.�$��8�[|�� k�#Yʤ�$�E�@���v�T!�`��4*v�#W(�ݵ(����Ŏ�:g3]��qUJ�FCC$�<])��:����n�pr�j�,wB��ꢸ��;g���qbD�8��.��J��a��ag���g��/�q}ߢ�voD[�2X`����;�S;�D�jީ#d�祕"�Y�f�͋'���V�@����-ǲ�Yʚ��v$i����x�3�I�R	a2����C>��~N�ђ���SCؙ�Y����A�فzo�_�r�� �&��1lY�@)F��ہr�ك{)�X��o6n����U��h�񺺴i�Δ��ۻ����Y^�=��NҁB¸�tb��C��I���f�->QO��������H��i��f(	 8��4�$�+=�rۢ��8��2�6"�~գ�o��R�����w���/>�B���G�D�j؟�|��G���eS������<��E�����g��)���A���yq��ow�ۇ�,p����O���˒��e���qn!YjY���R+Oj3'��)�E)��g�Ҳ�i�����8���?wa�Дۀ��[��7h�y18�Η�����K�=��lV$V�!�s�ގ��z採Ql��B�e|;��2Y)�]0�:h�rv�����> �l�ۚ�ݍ}�wo����P@��6
�b���b��8ot�?�.�d�l��ʐ@�Z1�q6�J��|�܂D���)y�E@E� )��1ʢJ���Tnڵ)������?I�033�w�d�ΑG�Q!���j�Tg��E��5G�B�H��a�D ǹ��<� ��$v�
�"��+�0�	��
�7I%�h�B�S��2@�x����AK���W~�|7�|~\������Mά?$�m�C�$|��Y�[�(�+[��XC5���]���9D�8N���c[���T�G������[3/��y�W�˯>CX���v��ˠ����N�`b�W��NmF�z6���2��@@e양v�a��QLM�����Nݩ`��"W��M,�Yjdz4��Q�������Mw�ŲI�1mr�V�Ivxܒa4����Ts ��j(� N�^���Z��t�֛�����p�h5�}������5��8�>�(�*�#�0��joU�E�Q~)Y@!V�+n�nX��W��	����I��n�w�7;� q�˅��3�ʅ;�o����᪫�u��)Q�"PI��0��\J���e9u׃튶��4!�燰��	�_�HJ�B`���@AM�9�1��Y.ZdK[Cv٬[�D��xE �ﺔ��3$|\Kj#��{�+�V��<T�FCi\&8���B��F�{�(w3�^a/7&<!��d�G���d���e&��A~t���'_m�=#c�F���^���%����|��
�K;Uڔ����C� -�M�>
�C5��u>�׶�?L�ټ��\9�+�-�>�P�@��B��#*yΚ��+
�~rl|X�\6�����8Jcvc����� <��: �`��yLx�;@�A���DF������*�k2�D�0��e�)�Zo_��$�$����*���tTHP�{]�Y6p����.0:ڜNö��7��$[���g
��b%��i"�W^4����)H�b+P~�D8E�j�W6���H�&XP˃`K�`�&��7Z��
mga�w8Jto�	�g�&^��o$�ֽ}�=�}NhC|"� ��l��ͮ�����)�̶5d�N�؜��ZK-�׿r�D�=��9��KQV�CX\e�"��1h��C�l���f�G��_�:5���%�Z�N�;&V��|���j�r �����hR�)�N�|�i)ۘ�~ˊ�L�aCz�>k{�;_����ěA��jR�����J`�ra�LN'��{�G���6�)���85Ú�,�Q̔�;R�L��v�<sם4�a����5��.�V��xU���p�+Uۄ�Z^���#�Ͻi�	r%l�1�#T�ʂ�<���V��?��b>��u�>,�������B~S��p�����=�w�a���x���A^-�c��YK[R��#�&�fϏD�Qy|%����&��>�aW�Ŭ��CV�� EIη�������%�VQ���.���\1P��I�&5�c��V�G%����A��X�k����WJ�:�)c¥�=@B���i��{oY3�qy�Ġ�F�b��G���o���)"i�ue>0vu�2����Y4��^��{�⌎I=o�q���K�b�s���2�E���Cr�c��#�/�ڬږL�ي;Ԫ� ;����Gb�.	1q�W���Ծ�Kӑl��_��a�޹Z��Q��w)��"�H
��? ����(�fN�v0��Yn�yCu-���#���I ̚�ŸǤ��f��̗�s0Y�o۫uB4���bk�Z���aL���g��t�	s�B�ώaZ2�
t�N�w��@�~�Dko����Y����~H�~d�N�m|���J����ڜ��Ìz���pq�9�h������0�j/�"PZG�5R��p_0��Xb����V;p�E
�rm��do��ï�i#�Lҙ4�NvLg`�ؘ\T�~�xDĀ�W�a�yA�t%��� ������f���ݵd
�SZT#,	���Oõ�Q���y}�݅��-�o�G��j�a�5N�>	�ZD�kl��[��&o����0bȮP�0S�-g�i��8"�/Oi���@��Ox\�]� :�R�O⊄��hh�����:����T�ڕaW������u֛rY��	nO K�E�
�J���qi5��8����k�i��� #p��6^��Y�X*R�r�A�z��DR�Z	�S�낛�G}����b�W�K�)�-��<�ov�Υ �U�u����>!�Χ��&��|����Q�0���F���K	{�X��ɏӄ�GΉ�h�5�����ڷr�-!ה��i���p����FpG����01��+P��z�����d�Rx�KZ	��2�G��|F�0�y����[�F��F-�IC}�8���E[�@`�>w?�j�q�,W���W�JJlV-T����ҭ��t.��k1rnY �Ҁ4�*��]5	؛�;^�S��ȯsW-w�%���#A��v����*u�m$tz�*nz���� x>���i��v�ψ�`Ϧ�X����	��=�h$-��u�.yE{�ߖjo���2�?��I,f�]$����Q�$������A[v-��s!�c���9��@�-�2�m�/�M���%�q�M�$S��A����\��[���|�YlA����R�ځa��D�TJ@��U�W�Z����:����r[�f��Z�>�u�����O:�
��X�ˎ�{z�r>�Ĕ�Bo-����C�H� �ԛx���J,&���@�O�A�]g���X�5f�Qܚ���d�/�0�:閃�f�>���t��̴��3��_]�v�=&)�!��f�r���3k���7��`�����4�)s�y��{QO�^$�R
0��-w�ػ��zdu�o�+�>��A�{�͠zj��>�`᡹������R��w��lT)@=�Not<���"�����oD�ťZ���b	��|�K�ϧ�����=�� /h%���K���|.��F ��Σ�;��֟~�V:Zi��8�Q��z�(����]���I�
dP7�5��"�d��l�Z����50���a�Wj����)�C*��s���*"-�Z�� =3o�f.q�L��E����LtðJư@�z�
BP�k4��%���W�M�x��?����)��%6v�m�\�m��$����W����k
P�O�R>��q,j� [D�Ow�N�j�@k��|���+��IL�Idt�>p�bS!J�{����?�]X�ٵ�G�d΃�̥�<�tR@��Ӏ�<0�=ʐ���܏-���v̭��,��������H�����"$�0z�/�xL��Q*2��|�4��ea���2�^]���T�床��C}�D�ɠ��W�]��N>q�������*Ԃ���q�pTGˠ��1�՞���c�v��jV�������kޗm�M�z@��+��(%���A���s>���#�Wi���@�g	���(�����V�"e,��u{�o_���^D�G�V��I	�{�X `X�v��M�҄?U������6���J�լi��7��x�a��jxl{��G&��~���Ym�r����	N�9�c0|r'�a��<J�!?cˬ QG�&�+�p䍭���z̏ :�qk]W��<��̏���d�zr�\hq>����od}�Q3����{TY��+����h&{<��U�TQ\g}T�O�p`&	�������/T�M$O�VsK<HQH��Nk��9��}=�R�����Cb��R~Ǐp�+��������-�&lȹr(��7P���'��b�,|}Y�޾z��j��P8�.��8��m�a%^�|��Vq�.�'W�~�I���wb���|���:���]��m><-�6c�,�2���@�L+���. ��#o�ٕ�W�¯��;��ϥ;��2�*���ptҙ1%��ATUCAC��Q�y>�/�B�s��j��k�F9�(�8��W_|������\��n�!c^+�IK�j�����oݘ`e{�;Yee��Ǌ�<��ooF���@aݙ��#��ɑ�gw�}ؚ�X��ä�L;��F
�U��X�*�޵;F��2i��S�t f��
�=�SG�%�^C̷݁�t��wv/�N"��k��m�Zq��U�^��fn�x�q@z���RR�9�ۻ�zs�B��#��!�u�������2>�X��o:�cS��Qbu���)��雎Eag�$fb��G���Q�%�8f���+���0�wR���
��]��5�n�_�{��������>s���}x��0U�W5)P��,R��`&���uPo����=>�*���p���y�>���w��zF����(N�d�����u�����_?�61xv� 78$:Bi�o:�^{�E���7]îϙ�#���qgQ�Ђq���F��M�����:x!���.��E��_)W' �;?Ę���X�;��H��N��U����V�i�:V+�2BOl���E"��J<��㓑�{�K{w:����u��Os`�OZ�N� ����'�S�H��(m�{���o�VR}J�q&5&��9���F�H�xM���f2&uйc�@�y����᳼Ic��h;;i�O���ሁR{J�!ޕ�(}^��sWx�O�v���,�.�5qϕ%��ߙп��o�{�]�G���Yqp�1W�K !������ d�J2Q�A��^��@h�e�0��7����q�ư�^�{�߂G.�>.��((a�.Ԥ8`�	D�	�Kbl����'ȩ @��t
�Q�?׃L��l~��n�����].O!��^�'���xM ��"}:ۭSG���>�
~"�\r@8[�_ۋyBjo^�\<�W^��# 
T�[�Wu\�[u����t�� ɵP�l'H��Qb-3��ٵ(a�Ʌs��$m`�%�x�{��ڬ>z@�}ß��Y�b3�������`)]����=�現9u �"�j���B"�����Obd�M�B�����q���Zp=�b�?��q�vf��Vۛ�١T�#gu;�	���%?o^��,�~.v�U�����{V�؅�ʰe$l�5i6��(�� ����/eq�ᯛ^'�zӖ:J���H����n�>@�����Hy�w^�6����I"�p���}J�v9t�2D��g�3���g����q��@F��y�0j��@@CB���&0A�l�k�鹨��o�z�ZU�� F�����Y�ﶓ���+��@���o����;�����PT�va�.Z�[Y�[�M���ir�=CR�c�H�^��G˲������Z�:^�SMG�ђ����eF!�U�̙��f{Rc_J�$�Y���"v�������آEk���� �[zO�	�{-����ߛf:ӄTr�\A��OZ=rB�V��Ǻ3DC�]��7W�Ie=�%�V��U���0�4���}Kk{x��4��TPVUb/�ә��T)��p�X�w��oPc��xJ�B3ΊƵv!Q
@o1,�Xu�:� ���_��Qjw��a�b��/Ɍ��EoǱȀ.��V�?+ӥpE�go����fY+I���o�����0S"�����o5�pF��3�5��H�n�F����0�|[&���5�.���M�74��[�x}ڜ�f#_t�׌-蹿�]y�"V�3�9z4����|���f��q�:PNy��h�;й\J��Ԓ��y�)P��?@�|'�c�eV���Q1DJ���MNP�0.���酏���XU�b�����ں��=p�{]�3O�D�涹1��/�k��'/�V��O��<m
��.��nS����o��1�π�"�{�~�����5��e���^��ؤ���*��a�)�UEr��I/{nc�RO �D#�P��7�tv�6�޾F���m�.ԙ(����� F�>8g��{,)��*����1�!���L����D}��ל+C,��D��$г��J�f���3���P���\ZB����R�ǜN��(۹�A ���U��,�ɢz;>��Q��\����4�m�ֹ�"ТiwвS1�/��#b>�[�o��o��$�d �_fx-!5-"
�VZ)��?.i^�05����)���#^�����v%iq,�!�Wg��D�Mt��DI��ȵ"�E�1�\��-w����4�K�	.n
f?nDփ�6V��?p������Z���[�f�i��#�"
{&�٦�I�-�ޥ:�[��|,n /����iX��j�7\!@|զT��H����!�H��������6-��+��#�o�W���8u�8�M���K�䊣��a��{�mnX��<0�cTS���GI��
D����sJ5���ڮTsAv�:k���8f�#y�!3���[X6�+�j	7:�� ,��� 1Ή"��ܭ�ˏfm�L޳�W����.f�	��.���n�t;{�[\��Q� �j��fa�PIRC�X��:=U�����KP����5��sQ/N�r3���"�p4	cK�?N�z �J����vy�J�r�Hk�O�>��R���5�*x��癉�z��
1��봉�˲m:A��\&=�}bS���`�m���]�?�KiN��;R=�˪o������F�f%�$C�4z(��%���V�����g�tY:��A�L�cP;� �Z���j���1��u�����p��M�[[hr��O�P?�(���)��Ps��~�ϜfT�Jh\pM�������1�Gq�,���#�d���NTux�J�ꥐ��C�A�_ !/�nW�*�[�ZEX}mdni��*Tp�<<2@��-�P�y-t�c�ul[	��+���1g�J݅}����%0�%
�p)���6�^�=~�˂������'��u^�I�� -���<&�����PPM��&���\� 笴	�+��S4�`{nc�r2"�@�}��Q7�W>�k���ۥhA��c�w���1�����#'�[j5d���8��cRR�-�y��\5 h�4���=ءXF�<��yBwP�^1z�=l��(�F_�������.��r�hΨ�|_�O���gE��S�2® ���O4�b�N��$�=��B�a�]"�U�<b´Յ��'s�;�/�)�Cg$`�DH���P���P�ķ�����qY� ü�p��./i�/�1�W%��	H�E���	�J߼�i�"�/q��[r��3O"s^Տ[�
�6�JTS{���W��R�x��d$�G�-bU'	4z��j�҉cxH:�w��#*�`)���O!䷛�;y898�,�@F3�O���"�YY����
RT�ڈ|�+zC����[��yā#l(�)＆��MH$�-Cz)��|};���l�*��{�Ȟ�"t�~>1xMUt���{�W\_�<[��$|Z'ā�m�t�c8t��A��Wy�0��q�B�G�,�d]�|�-����V��2��k�.zT}t�	��ӨL�vz�"�Q�� | 䖫��gk+7��w�����im ���� a��5��4�Uc�ny
��XS�\�5Jz���(��
���1��nT�l��!b����n��%��U�Ut�ZZ�ow,����	L��Z�X�Ֆ��; o��^�Xp6AA�l�5��XU͛zEH����^�������y��N�X�-��-æ/R	��&�m���u�����c���td�]��xvH�/�#�Rw���&f�|TQ
���F��.$ՂT|b�����D��"�d>��$���y��u����6��~g�6�]`(n�e��M`��-%�o=��g�����q'���Q&,�iU� �m���K#H�%�2���kCʝ��h#oYL�����i���j�O��ǂ��+:ԟh9&ͻj���<�4���ܭ���X�4������4���RCr�/I�]���1c7&�γ�-�Ć��Y���י�-��FI� ���척�X�KX�Ni�Q���.3�@N���J����wc4��)iz�/9Op2zI�n�t�+���v���~����A��U���{��+>RP�g�ƿ	�� vvD�}�"X���sx	l�)�!�^���8Ȓډ���h��Eܒ�`�gV�j���fZ;gIOK2tô���5��tz�������*�<�]~�i�f�B��@����ϰLigᘆ}5y�$hsՌ{��u�{z��H�����ni�\�����wD��=����	�u�*������/ �C6!��7��`�L;��墙���0�vޅ�@ ��ͳ���&t����b�j��g���PI+����a܃�&��̐u?��7��5
��J�1��>�S�L<�t�Ѭ%5^8���N��B���2�+E��U�p�5�.2��Fq9���D��{�qj����U���\@N�h���W�s��Quh8m4W@�R�6{% ��;��ċ�^��E��-�����t�x�%�-3���Y�w��L�/�O�$@����bw]�{��Q2=�74C�B��_�����ޒu�p��g�x�?�}^�>��v\]e:˵UO��O i��Z	,��xER]Vd��6ۓ�������'���+!$ ��AN���U(񡧕G���ص�X2X���L<9d4�_D��@��n����ƶk+_�5G^rU҉-5��`j�t�k�L���9ܴ���}��JS5�TS�[�;/{���z�K�l����{iΌɭ��*X�+��j�
�F �mz���3�R8�P�^��3:�z�T&lE���T:q
5WfW� ���W����%�D1�,{Ί�~��Z�G�~����`�M ��⪶�kX!y�������s[������P�es��(�I��aےPw�)a�B� �(���o�@�6�z��L�f4��Vr��e�di�N��s��[�"30�d��}V���]"ae�����h<?y[�̯�PØ_��Q��<���H�6�ef�+k���o��~���4�b1�)[���o��w2P`��+�m�a��j�)Q!�% �c��sC=J��-m�B���������,�ƴc7��9�b���ą�D����τ�&覉�]�fN� �X[��<?`�e��V:�v��r��]i�z�s&� A����e�щh��kS�%��e���~#NV���;W`�Z|c�S�,<^�
(��U,�XP�����@e��Xlt�����T��hq�ǚ��(��|�t�w|�#],�O���6Z v�f�?e�_�'.Y`^��@R�����l�鱒D�|0�>S��PX�p�c��
J��C�s.zr���0ǥ��yn����ͻ5��D�e�v�ŋ����aP��S9��WYj�H�#�Nؔ�W�q  L�@\˝��
�?7(�	�s-ر���Y����)��K�׍)3H;�%ޱF*
����D�x��G��%ES�.�	���/�Y�Fʍv�= �{^8[Lo	`�Zb}��SQ_�<Bo��?�cM� �Z>5$E|m�;�V����%�i��6;��i��ROn]�V������w2�gب�$XT)Zˡ^A9U9���\�D�e��̷)!��{4�p��JH����%W��j~>�Ϝ"&��?�94��)�B������ȑS�T�>��?��z�ȼ�C0�OU����m�����C��SD�߁��år��ە���N��}X�g��+��XJ���?�\�[f%��,H�G�$��>���B7\@Q��q�,�$�y�jRh����#KQ�a.������xe��G�+��Da��G����r�&vl��B_� ������(31���S�&���R��pL>r�ih�1��z?�ә�[�5�����⽢���]g�.H �+OY�pJv��[�rw.]�]��9��3�_���:���k��u2s���>b��g%Y;����7G��,��:hN�/�ܪjĵ-mW�X:
��tOz1�>yH|�ޤx�Թ��S�e�A�bR�(��P�	�*[ye�-$8ۖA��YaZI�ޟ"$�(���b����ӽ����G�B���>*�=��'M���6\��,Ċ�~�R������Pa��I����^R���6��{�=&x�h
O6�Q�`���-w�`EA�}�nӞ{�eP~5T!ҟ��!�n)�yө�)%*,]��'G$S'�������u���8�Uyi�Zif1֞}�!2��)�S@��?d=�
�����g�_BT
��{^Ĺo��B��A��D�/�":�:��;�H$�:�ݚ+hqs=�7*ʄ�kz��� �%�)���D�=%q��E� �Ͽ��2��6ѹ�զ'�"5�	�/ E���!̄Y�Y���$�����7����?�r�rg�P����Suk���	f_�\��ȧ���c��q lM:⣱r��3�MK� �dl���js���ҙU�r�p�-�H���r|T�J���!d��O&��D>�fK_c�!���%ↄW�=�l�@�:L^�I�#��R|d��-h���$fVL� ~�\H�V~��J��`Q�����"91/��C��UO� AE��Iw[It%��H�l�1m��UeȺ�a�\�hB8x-U�^�'eʕB"����\-!��@f񼯿�~Q����p�ln��k�{+����ien��-�{���(Bu��,8�3!���������W?CpR���R�Tjk�g8����,Uk�ʌ�@��7��ea�"v�䛇�W�}��|�FA��.����Y�o��5���[t��?������~�*Z�&ɇ�2+@v�ĉ�� ��{3~���X&�$j"���sE��s)$껝!�ח��P�8�ҤZ����C$<.�`�Ul�:�z��Ƭ��r��PGKN��f䱒u�	���P��y	uX�A�fE/F�ātt+�#�+�ppB/rB}�k�8y��/w#W'����7�Ʈ��'[
1s��3�7_�N��.����T�����m�L-@����4A��:rrK�^rT ���/�o~���?�$H#�N����>Ց�e����ޯ���,�D����X���*\�}<��O�d�u����&�X҆��M��z� ��nj�D��~:��ؖ+���'�v��F�����-���h��	:�>Yd~+rc��뤓A��V����*�)��hggT���I)�^]G3ן��D����a�H�9����8���K���46�6����FD{��<�)���Q��> 9W��7쀚�� �@���"���kf%T=���ݏT����_	қ$���o h��bsn�X�ARP�a7/��"�h��R
����W��zJ� F�t]���1���TG2��d��R~�\�r5g�E$�#�N�z�4W>����s�0�(���'�P�2���4	�����4&yӰVci&���*ŕ��X�0|t��F��@�׭e�ig)M'��Ʃ���lB��b��v��t�w�z%�ЙLz�����w3��U�޹ ��&V�-���
�L��<��~��P�lQmT��j��wӽ�����0��gc�ż�h�Ox�`�v 瀒E�{��Q<w���P9R�<uk�V�q���_�Rb���~�-���D��D$$"oQ����;s5�j���Qi1�ʹ�$�z��G*��˩��i��
!�ĸ�`��8_Xtvv���H"LVhh�qx5��Py�wna}���n��I�ls3?���XX��!C�'��Sryp���9�v�܃c��
��_�9@T��\�15�:�W�}U/
� �G���S����(�&{#*���(K�b_��ԘmR{��Q�WşI��V��q1����16��*���<�Zs�1w��&��8�L�D-�u1����/l�/���D�iނ_�,�,��� �9�E��Ʊe�XUU�lu(��)�j���V[��}����]pO>7����:kGv��r:fi�>��Z?�����N�mȐ��nu����4e�^ê���]�(;	�����\I�a�d�������WK�ͥU6w���\i�Q������d��n͢�&���H�����������G�:ί>^m�+%�ˍD��"����$(����~$�v�����c2�;P�x��l�f su�66+����|ԯj�Qxx9�7��X�Hދ�2i��(� ���ꪻ�
�{1���B�"!�W�_[Um��AU��H 	9�D���v�{�[�z�B9:�I#y}�1Q�L�x�Bz~12�{LR��\��L����!o��1(k���#�A+�D?I�ͭ@��������m�r�K�2]�9��凿 6�9��Z���	�fd X�c�Z,t�an�uA�����]���������;{�W�Iґ]T�Ym�ِy&��c$u�-�{ד#n}e �>���!�򏋒�(���k�<�x=v��Uq�w�Q���U��=���.�o�O� ���o*����-�R[���I<dfɮ�Ip$�Η�ϳ�'G:���D��bf"u���>`�'r�q6mx5� �+������sT��˅�1���ý�6�Nª��U2�n�+�b�3܌e0�%�KgM���Y�pՈ��}��j{t��dr�{��n�@�Ipy��F���\¢TAu5�;!���_�ѶB߰x��e����4�9��u�m)d��~֪S���Rz�wᎾ�uRpc�ܽ�c�"����X�TƆ��n^����A�ݪ�R��C��}�L��Ajcv4�:8����U�+�V����eyZ��O"��YguD}5�t{�B�G�B�+s�%2�r�[�=�k�+h6\\l>j�;>���q\�^�Z���׃@?�*2�JN?��ЧB>,���$Ψ��^i�E�������(L�J�	]A���c�U>
�eB��%9����U"O%� �V�>Yy���� [�ZRk���*?������>�rL>X3b�s�P���:ü}D.�K��ku�8XPHu�\���2y�O��yJ4��j�CBICCW���qq�{������J��*{�{�"e$�[�DR)Z�kq�Ɯ"�����d^���(��Xe7���ы���ʃ��g�.�[��P�;�ݻ*/p��a[j:b�sR1;lh{'�Jꊏk���HcӾ�\�b�5	�-|Q�K�����8��2�.%v��2�_���Ы���g
`�����ѢO�q��5|4!� 1��	;^�A�)����7�R�e�'*�{�աv�|nVs�3�LӁ��$ct}�� ���ap��Ƶ�.�z����糉,�h�r.G�}j��lV�������2P]J�w��밹ё zBC�JeJwFt����-�\�2����9^�x��V�,�2�š3�2#��D@Ʉ� ���j�&f<߼a[�ݍ�&,{��W;z�@��Z������H�i9�P����?�����|�������jM@E6���:|8�S��m�`?�7�e&#դPp�P`I�l.����>ezj^x����b�7��ęR�l�����C����+��4/3�����U�@�X�wCY0W�����O�X~I��ط��&�O�,�їĲ��&���nLҤ1�Gth H	R,����8������ �,h� �y0UؿǺ?�������Z�35�ɋ��Vӓ�߿7�<�g*4p� ��h�o%(Z�$�A��n|�PE?���,V���&P��=�����g覍8�>R��ɨ8�����Ҋ1nQté���t`�e��	+����M�=3�E'-�.7�-�%���W��ܕ�Cn'�ʌ@�#w�^	���o�PS�&u}z����	QG���I.�:�%�ch`0œ'-��h2& "�:���]�5�p�?oN�֏45�FC���j����0��Bg%OQ���6lp�>��<Xu$P#�%�w�)�]s����h#��l�v�_.�8��W0K�/?���c���#\D�+��/vt�29؆�#�N|>+~7Y\"��9�kns��d@��AqA>+���=��_6`�b��A�F��g%���+���� ��,�Z�V,QRْn|��b�D|���7An��i����Ot��j3��0R{��xӾtJ@(��v�a�@����i�=$Ŕ�j�_�Dw��-h$߫�\�8��>�TA�.�I����CN�L�.�GG�����k�v�A�ѯzj4�Ǩ���B��eڌyC�U��bޥ�{��6�`���F���w�h�T'�r�P钮��D�7�N�ŷՑ�E�.CW#����Է��t�н�b�VkB:_PC���op�9���hɫ΄e��V��y�:�^#|/]���i� �u
�j�D����&0EƦ��il��In����@�m��/�1�ϑ"��}��2�@&N��vq��$��x>ߖ�j*�	�)dv�!�.dV��l�8 �X�B4�F�i7��^R;��gH��ͺL1�S�����0Do�(��Ai }6�4��\���W�9}Lc�J]~P���owp[����'a�����Vs�fq�������ϼ(��ئ�mI���I䳀N(���x#ER� ba�6��^s5�ykB�u���ß|�
�S8��f��q�N�QfR�v��������=�湷u�;Bl�q1��#�s-�k��j^��g��F��@�s@ ���a�8���2@�ʾ2���貈z_�ԧ�b��[�c��*
��-�u[�*���^�Ф�B��XMX{�u�m�F��q�T�'����07�L
��x��{\����fT���*��a���"��2�^�� j3,vL~m���z'Z`��	��q�χxV������K�J�S���Ӷ6O��"و����,���xԛ/l����'R��V�o��6�[ۥ���Zʹm*�#�r.�}�i��C�4t�.j9�K��f�o��(��鱁�>�y�4+��7��E��v8�͚��9��L#���|�r8ZR�b�,� �L���~L��)(
��k}Ҡ�G���b=u p�.�0�X�V}�Ѩ�ozx���S~d��2��I�D�F^~����C�+N:�B�F�1Y�q+:{��=�_�}a�@�����WɊ��1k<�<S�뢃���|=���Sی/�̚6���%оe����n�������<����c$'%�Lӛ����o��AC�,���:w�97(�)�,�ù3V�,�2c�4;}l����w� �f?O_>��L^w ��M� B����?� ��KʨF�)ɗ�Q6�L��D�0�>�Y���FL�NO�a��Z�ia.(y�&�H�$�y��$��_�k����Ƹ0����KS S	m�p���!\�z��|���^��M�˾9`~2���V�/MD�u�;�F'#��1{�S�N���6��'�ۚ[@ۼ���K~��U~ �~�^w�"�<��D�y�b/����`q&��z�W0�����a�ɵ�Ƒ�=�?�ў�L�%F�}�P�x��u�F�~\=����	)�+�{QI/w�Ros��-[޹��s���:.?�Q�vw{��|k��]��V��E����O�z�ߛ�,��Sa{5܏,@�3���4wcY-4�D}�M�,��(M:?���ìT��QIO��/ܬ�]�~] �AԌ���
۷X6B��¥-���H�n���S����.ΪU�{�+��o'����*/Rd�<R�| �A5{��5����I��[M��&�㧒ڭ���<����#A	P�W`�]/��ީ�K���K�	���:�F+����ʱ�H����h
ֿ��T����9'��ܮ<�u�#�#֨��Q��ME��Z*��A�e�����@����C�mO�\�EO3�s	l�M����>Յ���F��<�#s� ��`��>/�����E����a��m%]p�ٝ��5�+�ާ�<�����Y(,�v`�*�E���o�U6|`US���T(�� �ND�s=�Z<�Rï��&�4��P�����^fi��g]\[�lx\�A���WE�_;#F�֓����^S���?���h�z��2�'��m���Mr�F��P��gñ&������թL#�f(<�%����k����9�<���ط��7�Ck߆ru���^�nIb|Uɏ���.�d٥4�X�p�	c���ar���T�Ba��#��Mg�Q��waUMl�����2Ct�E=�~v%V�O� ��TET�zZ<Ȕ-�#U��� iL����[e"�7d�"�kM%	�G9���B)���/���g6��Sj;Ej�o�U9�����zq���0�����%%a#�1��^���N�K �̲�v�n�l���H���N.-��h5�dþZ�گ^fr�����u߰�I�&!�L�u4�3(��ꌲU���k9S��D�ԐQ��ɣ���3�T��{C��+#T���� �Â���zCض���mU��m����ǙV�?]�ɻC���G�S��Df�U���{��f��S�+#,�Ǎ��)cwں�؏��Aw���L��P�g��Ԡ< �x$���e�W�3�	G�r����y�:"��ƈE�G��O�%,��:i���(Y�]��3I/R�����͌D�������/˴�W������9�ke�4��!�&`(oA�\ԁ��1�:ee,��`��sE�[+P�5i�����b������i�R7�n�^��ҿ=4�e�����KEA_��?�C���M��W�^B��B~.��#�ՒY�Hގ���!@qm�:*���
[x�Wh\��q��j�F�r�	��N��)��UWl4�^�>zB���@���d�%;�8q~�ՈL�ȉ�b��^R`�7�}�Ԉ���J���E��Ћ���O��S�ʙP��2�r�wpV�z�,=_G�}ϣ�����5ˏ���_�7x��bQ������d�6�S��n��|L�͖�_!h"�ˮ�~�=���r���mn�=-��t���t��	�ب�����I�5��	�����c�wJ�X�ߝ���Qy���i_P�Ŏ%F۶��(*�xB���0���\C�@N�rB΁D�R�B�wv;������@� �1�3Z5���A�����p�躚�Q0�����ɔ{�\�9?=���3��-K��m���k��aE��m��+�����#�p�ES5��0�_w`�o��뒡x�]F.
����Nm��kA��ݖ���ᣕ��E���W/�$SĔ�&*0�5)�2����C���d���-�-HO����̫s?���Bx.Ƹ4|�N��=�Ē��!!z@��Qv�I�y�� ��q��`��R�"�l"�ң逥�mg�Uo�_5�툛���3W�/煜���Yy=g=�:"}p���';�&nQ�K_t���j�iP�y��m��T������r!-B��Xz�y���O�e�95;�jIu85g�jT�h�gh��ۼ聳DGg�.#`
5��������
����.��'[�;Z^���~�{m�Mu��tB1����uqh������4h������,3����N���<9��#q댡V'�jP�d8g��k2����!�L�h��̔������?����3,(~��C���P3�;��ò	Q�z���M�n-/H���W=����>u�X%�i���,��ȩ~>/' ����R���~������`C�|�K�k���G�9�:�YY�Ab$�t�-"!�9��׬A�����q�SM���&_�lA�V�k����X!�w�Jo�/�QqM�@j��#�EW6��ŐQ�춛p���Y W�Wɚz卵��q$�X�td�ͣ�3��Ԩ�ƽ�O�\����Zۋ������qb�ݣN\���.���@S�b5�9_%��V��=�ݮ'5\�C<л ha*��A0ۦ v�ĞYJ����<� .e> �`�6'#���+��R���T���@n�t�L�6�_��'�T��JҚ����$DE�MYZ���c�@�axxxd��n�|�^�oU�c��oZj����7Y���m8�TGO�U�=
�2d��g��p����W�R�,��*Z��v�K�L{@ݙ�O1*�/ȩ��B��"A߯�T�UI�~l�ft�{������x`(��ⅵ "��U�k�,�%�P�A�ҫ`xZ땏,�4
>��Uy�q�~��&�B^��?ܟ!Mߟ�C��Y�:8�e�2%@b��)��bz�NzR��D��9��"��="�FG�>�G��CE̱s��]���y)����z��
Ŝ|�(	�Us1ӕW��f����#���s�ٷ���d�i�_�U��C�9;�p�|d����E�r�G5�Ϡ";����YE�^* ���G�	�@�Kן��2��R�⩯� ��円/EЇfDi�����Bܭ��&ro��Hc�8�R�)`U1��w��	e�(�rn�@�~c:,_nbT���]�a�'�_M[rp���i���Y�B��+B��#я��+ղ����<��]�[�0��d �5�P�1���3⦮��U0X�����jNc.�2��Oǳ�p{�4�� �N)�	���#�x;�r��]@bC �c��[R�)]�����*����*���@3���Q�퓛X��� ;p2⻿{����{�w5�.���O�a?�7*��Pxs�*�c}�;x%<�Ji����� ݙ�']F�v�ǉ:`$Q�
[���'��a��wmM�NA)�Y����4b����������<�hI�O㒾�p�Ϋ�ܤ �*��<��k?����gBKc��9�o7���[شAJf�!�7X]~Y̳�q�����s	�D���.���݈�%��iS��y�C!w4	,ەtG+���U�6hxZ��R'��$�����|�Q��U(\���n@�D2�N}������-^N�Ѫ��5\�h;j��Gcg�L����Cy����,�M�� ��#�Y5�I�[�;#+G�R�T����U��賦���i���<i�Q O���Ȗ��ڵ*��v_��W�T�t@jj;��|�!#�Hajf��a�`�b;����!e�b��N�k��h�ʗ{�Kb�(K"���A*��O�D���텲na	��C��1>��!a�( ���n�c�����XK��a%�9q��堯#�zs.w	�9��JBC ]됹���@�3��QD�䉉�<�l[����Qd�Ȅn���!ҕ�~��N�C$z���j��"zn���^��������ȩ2��`U����{���w
�:2��2o��3%Ӝ�0��~�H��K �������;2]�|Հ%��C	YiڇŅWH�Ɍ���6F�+���=V_�����
}'�G�l�I�0���D\+�����N=_�<�t�����H��Ǟ}�X���X��@D ���a�8ܞ���(It�6u�&�sek��S�u�B�yA�;w�̥��Xɘ�(r��=�Qj��5���6,����]�i���qH�"bc�4rn�"K����ˀ���Y�缒���o�]��
&'���A|t��T|���
�4��ȑ��3د���+Q��>@xm�����yZ�"�:�Sm�:����*"K��&�MB����0P�X�j2SBm꺀Y~1��F*�Q���}�/�'��gW�ev��9Mvl�g�������:��,����xg�H]��_�,9 ��!U���qP��ߜ�����ȹ%ma`'�E���F��u�V�:XyBd�^-�[dF�^�l$>w�������י������J�4	!i����]"�^�{����ݻ+��%À`��Ĉ����j�']�x���-3y�ދ��`�2nmLN���CL�������[r��J�#o@���4��G�D/0��K{��V��v*����U�|S̛�[�	��I�J�z�xXrH��Š�l�A��1��q������YV��f�mBhD�V�I���h�"��>m~��5�1�&C��%��k`7�GY>�Ժ�x�q?,�ҧ9PHo��V�&F9[�!E61�f��[���g���?�q��D�^2�>�?�;q��;�ak�v�P4s�ك�!�kyk
�&/���px�x�HI<{��2��Ո��8M~.,?M��`7U�X����2te�{���H3�\�|75�=�Q/G�����k�ݢ�`n4�*q�J���ڽY@�B0F��`��ĭ�I[	���vTj/jr����o��X�*��S|l*j3�*����@@�2᧋N�Z�g��-��Qi�$���o?�A%J�e��EX�E��z��ȡ)懐��v�^�6d�3�2z������1�|5t��~�\NV��\D8f�?ɲ�Y���L��h���vGHc7�wX,ƾ���B�S��$$@@��s�~��,h�3�Y�;"�s6\�k`��J:7ՠb�3�3��ϐ�W!W ��-\�;�`�a��ٶ ������̻���"*V�|	�`�bB0����0k�`'��A��X!<�.co�S^��$�)���"��lT�������fh^s��	�U�P
y�.R�g�~��|�%f�̫}�%E�x�X�y4y2��T�T//��Mf8������UI#p9�A��פ��R�<N��v�&b[� ���0~{�4Y:hGV0(�
,�6fW�\��o2�{���T�<뢤\�WCq郏 8tF�jY�=Ol�ߙv��;�0�b�f��(N�������@t��)�ӥ�gb�l���d;"�Z�1�81�MbAK�t���
u��*�Q������n.'g|�����bZ<,��q��-�:����t<��^�^=���
��W+��H-v�{�عJj]:��D��.�KKዒs�VD~m��������8�V�ƏT$(�7	n�.�i��� fns� ������u�Qh-hЛ�~J��(���q�A��f��V�3��>1���H�^��
�e~�����Ow��ލ�E�!)�I������\H���R*1���A �?!U��W$=F��ր�-��1'�`� ��:A��QvfW5���b=�  {�:CA8�Ԭ��8\��+U)L��z~v����ۻV��G�ې��+���l7��+�\�Rl Y��d1!�O����>��̳hM�՟S
�h����(�6���η%��4�ҽ�ߛG��++�Gd�;dv�@�ݏk���;�����v�$�dE���\��������#����r��O��>��*8m+%5�2eﭑ�.�[lzzq�S��R(-��as��x�4���O��]Ԃ�Q!7ej�S�mX(�'M#��*f���t�فS�4Ft��G�-���Y�Ŧ��_F��T��y�sqWI���/�qd�֡4��|�tqm~���S���F�?4�=��������5�S����|�c�P/�ywp�Vfysg�ݤ�r��~���?��u�dp��;�u]���kJ�h�!�Ҭd!>�hM}����AN��{��h �_(����P;ܑ����-���	U?0��h��nժ��Y�dd�S8RT�����`>�"�Y�[j�'(|K�K���Y>�&���\`/�m�$2���ݕ�m$Ά"����P0W*Xk=LHE'RT����)GA��o�!m0Y��u'�����voz[�<�����)�_�jt@��V���P}����hokY���M2�`O*�e��9�0�
`>7��=�_�$9�=�E�O6#-?�X�.�<%n�e�$���vY�\�QVA-m�êq����J�:���3� J+?e��`�iJ��J<��}I���Z���ȟ��-^峏�c�X��'>�������׋���ƵZ�g����GoL44��ڈ5ӑ���9�х" ��xq��qk�F�7L<(��A^ްW$W��(�M�A�g_�fI�L�8u��AiՖ��C퍘F��ylM�Ѵ��L�V�%��S�i+?$ϽL)���p�^n���ܹ\X[|�|�T�Dk$B�j�gs��{���T�B.뚤	`�"���vH#� (���I�Z=��(r[���L�:~������90$@����&\h��!��0�8:�N���J�Kf�yy�~�Ҿm T�9�>
�Q��C�9��!��V�~)4�X@�д�0��rF8�#}���	1�u>F�)x3����we#C�WvV7�Q��']S�"AEy�$��D�#�VsN�u��Z ��]�"nN��ǐB�ً{��u����,�Ro��[+����YU���?^u¢F4�4���]=p�$�ZQv��a^4�ߦ?�N[�?SV-�W���5�1����s`�ko����V���� ��˙��V�c�׮����z�z�2�= #�`���(-��:�v��H|e�,K_�����x�ט����D�_'2�֭��?��!�cu�O��Ki^�b�@���ٴ&���.�%�k'qT��wi/�	��j68l.Q�bL��D�����
n�Vy�5�(�3�s.YO�.{����]!{"9��45�"�����*�p-��͹=����τ���u��p2�+Su��C<m��Lt?Y��t�㛊����E�I�5C�;^w���oF@��G�ۭ5��+`J��B�U��v�	��%�X�*�V,����bgQpsnscJ\���b�L� @�hD@�=#U��Z'+���\dK.g�Ik'��̫7�C �yb�σ�;������Mn����4=�k�����i�SD�@3/��v5��Y��=���~С�����ޑ?K�A�4��~����S����4����z�d
�p�W��d/�i�O�ʦqm��𖦏�T
�D��+xB(�B�8pt�@�1�H�{�,�M����-W&��b�ĩ3˅������:YJ�)����>j��
*&_؏i�f��tOieNA0K*�:�$�	�����?^�D���I�E�3���Ǹ�R�8�5{b�vuM��� e~�ι�P�w�ź�M���Gp�mY�ɋ�X��8`���G���
]1r佰,(聦 ��׬}%!����g�3A����Ň.r&�G����� (��u���J
��B1�<+�Y#y�����y������ncl��V�&6T \��2��`�N�z�ME������E9+҄g`gxɺ/���Ok�8�֚���_��,+��B���X2v�B3'����'	�c{U���� �N[���@A�=���=����YPT��$�@�ve-9����Q>�.�|��=�7?��oH�3ֿ�~ܧ�mW
�i����Xկv���}b�^m׃��f�f貕�d�tp$�k������r�0H�mSL���yd�NK���!߲Կ�>wW�.P�|�0�y�F�UeE�3��gl9���s�n��'� ��_�+s�״Cl���Z='�ccRp�f��	��K���I��?>f�S(#�Q�y�T#���b�2|����&�������h+��>���"$,p�ER(��;�	� ����oK�ƃϽ����!�!CV���1���Ҧ�
�cCdØ2r ���\�����ԟ,7��2�4��&�p���������҄�{�j4Y��.�ۄaɮ�Zb܉Bx�%c��W�S�8�iLW�F��� �F&��l�j�
�tb;�kP�Yx%�W|M�������n>A�T����ļ�T��W����7�t��:X�������x{_Re��<���k���ΉoĎ��g5�}i�Z�CX�Vm �(�=k����$:�����s��GfUg(��,Bu�yOw�K:M��x�#�����)�Bc�]���uF�� ���׊�[�`cy<K�hi,#=�{;}����)g`�0Wud�o�xX��5�P���A=���㤩h�u��m �D���#�K߱�����*/KT]�Ҩ�S�*����f�.�.c���,~��g;�Fǆ,y`Q�!z�s�t�kyK$�ɧ��+�G:r
m"�G�l�i��(f�q�P!ѯ�Я7R�<pd���/J��������_�N��&NW�,�D��Э��8f��ב��#���m4io9����:N�B�9���)�Ɩs��,�y�$R�A���Ĩ.����q�L�|���~�+�r�v��R��������ڟ�_Jj���q�ga��N���ȧJ�Jl���#������F4z>�⎱ZK�+Vp��Af�w�R�n����]9�^�'�`�	� �t��:�s������&u�}��k8=?��~���O"
Τ�C��q.��W�;���nx��I�+�k�{����	f:xd�o��K��Oi�Y�
ޗML�O��s$�	�g����(���_;�'� �=���^�0��3s�Y��P�z3#���3q[O���[���©L,�J:�g]F:�,5����B�)�����2��C��SC:�P�6�M��}��B�Z���+��ZE�n�B��"#U�F�uJ�1q�D�A^P^f�!֟%
��:s�en>(��Ġ����������v���w�Q',ܸL�d
���|MN�k қ���B8h;�ٺ�"ݺ�zo4
�4q�ϸʅ��ZK ��Q�,v��Ně�mUE{�v��4{�K���ط��s��r:��80����%&&����C� ���gG�&�FC����r�v��'�W�����]���9� ��K6��Ə���A2�%�����P�f���-o��eM��;��9��lp�>�K�R�;�!�~R��d�� $���.��<��H� ��r�g�2̀�03C�Z���&v (��_S�%��9�5�,�x��ΐG�����3>ꋚ��s' ����+��VT�y9�O��E���LF];nkZMV.�w&nyy��XY�.6R^<fCfB/�,��Hh���h<]V�WY2r�t[��R�%R;�(2��6f�+�;f��}(q<�����W���M�b�+�1�,�M�ڔH�Q2�S�$0 ��� ^�z��e����wF�+��p�p�ɍ�.�dE~�&�ݠӝ`G�ab�����k�r���V5Ubs�9��b�_��ס'��.��dHI�]ڵ-� 0�cG���Z��:>��2 	w[��T�Dd��x���b��<�\mC�W(�{W�qt�w�rF\�������4?��2�I�Q����(�\�2���v"��h�x7(B���{�)�i1��5�>zZ?��ݩr+o|! W�O���d�����/#	{w��!�� ��@&��[�;y4}{�qO~��I|�D�Os��?N�q(�s�#�A�-%h�aR2���"�N��������lZ�i�4�ʠև�yәU�y�]�]�na;h;�F_�����x0^+D��F�(F��r���T{�}�i:�e�r�����Q�k��kk�tg��J��)d�g���*��V�E�r�� H�$���� }�̓�&���r�+�:{��C֦<��X!�z�4]^Fџ6�����b��
��k*.�ԍ�p�^���Q��Fe'F�I�r�l9�Kt/�X֏�էO��>��Ck�US�,Հ�ֱ�-�!N-����]���-�W�:�X�঻x�	�Q�G�mM���K����.����<,eO}��>U���͋6xs!��YZ��ySJ���Ε8뀙�����X~γ'�}f�7�p��^�+#��������}.<1�I��B�������<�yx��sp��^����
k^��_%U�|޳�*������O�@uW�������x����lT�K5w/����_�254Q�=�dN��^R�vi.i�������f�Vp�q��?���m]V�?��pZ�oE{�ᘃ<��;R-�q}w,+���3��BC3屺=�ǁ�e ��o��T��(]N��a�Ss������7buI��SQ9 ���;�>=Eh�7(���tZ���7���h���D;؏��^W����S?�����yV8��<V�H0�"Fj���bvvy,�`Fw8���=(BC��X=<Ӧ�%(D[����1�x���}7}�|�T96�
�#���h�B��d�{ˉ�*�%��N�S#v��E�`t1����u���A��֢��p�]Jx�U"u���i�Zb�:or�Oߣ�=~凙�@�!%���T�m�J���v��w&����ʛ&��f��Qz�v�ٞ�/��px�C̽�'q<@@l)x�А���a�=�~Yf�?�QH��^_���Q���ªA�`J�ϰ�ũ��&�K��UmU[^Ԁ)[���Z�.3�ZZ>�]R��"*�/�����pZ�+N>c�V��(F�s��0�UvJ�E/߰��-qA�)��ā�y ҅�Ϗ�K���O�9a�o/h$��l�).-u1H�9�
�fgo 6��G�􉐴'�H=�_p�����8���t%:D��jp���4;&o6�i�iM�.����=�h�z�'��I�)��D����9N�Pؐ�ֆS�]~�e�W���7�V�4�տ��}�X�2<�#B��x�aԴ�G2a�������ҪA�Ɇ��-q�g�/D��牮��~���iߏ����#���ɾ�hu�w#Z�;4X�%Et zhcul��������E�%�c8G:����&*涑�?.�Y��**�c�b����B�۠a��Bo���E0���x�H�r� f�
(��%.�p���K�*ߎ�w7u3ϵ�i.C�rP�;a���x�H�����(��砷KFn�Y�|Ǯ �]�Y7��;/�e'�� ;�#��I?�����7�D��%��L�� NN�����Hu����Z 4��][�����g�ztUJ�ׯ'�3_���vC�5N8c[^���bW�Q�oBrE�h� 
G�=�MO��7@�>�S!�C�����M�W��_V:e�Gx�ܩ��/��m���_����`��7�jY,z�^�ʷ������e��u
1����Y���x�tFӂӮBt��Kg*x�z�bY<���A]�ˎ=���{슊xN2���v��v�&�T/7��4�j�<U\�D��J�J]-q@��HA)�_�&ނ�fK�^����J% �����D�G(�w{$��\��)�8U��oL�)A5п��4^�PbVO#�O^�.��.-j��7��X�A��r]LNeg	(W��t�{���� Ӗ������R/�����qީE=��6D�¶�$ߢұK��������1��Q�c6MB鹆��Fy�]��C�Dr��O�PU͠�=#c�NS�a�-��i�<�(j��j��ԋ��S�������������A�\�	����%�����V1��]i��"��t�)Wߛ���aѬ�r��>�x�'���-F�1s$eaw���/@o��(���J�-o�sj�$�57G,�_�t�Hg�Z�ջ9�֝�z���=	���>�B+�}�A3�p�J����t�'
I�8x��5bI抒S�t��y_��%���>Qڰ��W����-{ާ'����krī�ny��=��QϧhC2h�ֶ׆,&ۯl��Y�%׳dr9+ғ���Cy,�K�aj��3�ba��])�v��]A;S�m呆�V��ON��ק���S�Q ���ҁŪu/c�ͭ��$?ۖp�����	] ԍ~o����rX󺑧	G{R{B��#�*׶H@U�9[hAt	ـ�9e�� F�����&�����]�΀�@ك_�ÿȉa8���R�GW=p����Q���mx���1�R��O����X���ް�I�-�֍����"��2x!��V�zrq�Lp�ʣ������o,ָ�_]`��~�!�}� =�dm|7Დ���u��y]��	�����4~ ,˽S�Խ���h�(t�9�T��)��k�t[��HlSMS�<m�k\�g���Ĕ��QjS�N=���f�?{1D��c4�g!1�J6��."]�|P���5�}(��h
�.�
�#���UpTJc�3��Jؐl&Rv֎m).?�;njtVJ�jP_J�8qL��b�WiYf��t8I�q�F(��C��Ώ����R���|��u�UQÚ,�_uQ�cz>�6Z�X��t>�ɡo�PeV��C,߲�M`T��3RxI�I��]0�rIK�*�Pu}_�b-o�o{����(��En�`�-
��Q��y���*h���V��.=�Lkߒ�m~*�w���J_PjT�7�lA��f�Я����o�l�ê�(�9����%�����j1�mv`vjt�N�֭5�.�/��<�8P%[)Y�W�.H��4%���C���GfVO�f�to{���Jɠ�j�Ʀ\m��٧�L�d���E>��D(�b���B��2�A��k��0�����|��.Uk����͏0�J�C#��%�7�	�B機0Ճc��Y?��e��e��a��m�e7��n�XsԚ-?1B�~��?(��~I����n7����=�|��f�O�b�~tK
�-�em)=+±wK�� �]�uQ%�
�a]���-S��J�`OW�J,��uy�K+���� ���~ܺբ�����6_F�����<.���p���QS��K��X�^��آpq'-�7#�����������DK�~u�ұ��Rr6�Nm),�#�^�:�ѻp�#��t$�@���Rd�~!�T�@�����[�-�5�,~V�:|���k�&A�����)�3"Nn�L��T+�����Q^�
X��çصJg�*����'o�M�Le�!�M��tH�%N�xC���J�f���Cf������5��8���1�ft#d6��l	����j��z�Rs�k��Vz5Y�~g>���[cڨ����@E�x�SK�w�X(�fo����۟�!���R�<C+�ppv<�wQ�xe�[�L�N���~�g��y=�ī`���>y_�:a��@�m��^?z$�q�2Y����J�h�9m�y
Q7�Ҏ���r��P7�w��;3�}e�%�8�To5}� i������ؒ���w��j||�Bۘ>������x���(��ؽ��f��Jo*��>������Rؓ�˟�/��c�t�-����Ԙ�6(�d?+�=��л�D�|F;|cR&����nF��c��?&�K�bT�QB�uޓY�5c�k���C���N���[tG��!Q�1��P@(�DL�g\����b�p�� h�Y�##��X���x΍��z*D,@]���g;3\v��!�]I��%��ֽfF���o�g�l~<_�\"��4C=3_���w@�Б Œ�`���빮���p�$T񄪠��4���`� ����ɧ���s��.v���� `������f9��s)���E�A��'�ԴV���t���	��2��; T��J������$�h6��2$�9��,�������ۑ��6b��o�hh,���c�k�ڞ|m-��|W��D3�$R95lׇ ��7�ꆄ��v~/��Na�FĖ>��W�`����Afx��^�m�띣�����6�m��|^]�R ��~�~����#�Z�G�ē����xq�lʀ���'8NC�r�]�y)Ao�Y)}�]�����M�c����������t�'cGA�[pU�o,�����`��SM�X�dh��H�Z�q��]�z�@G���Y�<ե`��^�WrO���ԟ��OX���yF���}��-���M|��v$��MpM����Yyj8��܈���^0̪I��o2���!�_܅�dF��L��oь�k�x�*�S���Ž3�S�RL�)�W`K:\���l5��M�s��>T*m�Bĉ�&�rqv�����t����=�2V�Y�E��%�{ǵˋ�m}Zeӎ]>� ^S��}������><�3ZwP���0�I������zy��?��bK��D��Wh���۩�����Ú�<�2���:�G(�[w�v�`�Ð$e1�ŔXiWlΟ&d�����m���b.#�?6�A@�1����x
@���J�c�nqWڤ0h�h�=�B��xFF�K���J�z{I�"j��~3�B!��� E����F>	�1���
�`,�}��u�__��s2L� 1Wo�B⩩��Y��	��_2�%������;��957ݹnQ���ew<��Qh�C?��韂���[�%&>�Pre8ιC�y�oė~�SB}���.�]Z���էq�8��M5]&]�����Tj�e��"�H���{�>/;�uD��Z�}���_b���}�'�)�1�l��D8�����>�΂C�B��ŗmêM���֛+E�mfo�� c��&�({���`�U"r�ft;T���^���!X��� ܆n�T��d���L�#7�5C~v�R��04z����(�۔�㖯���]�ŭ=$!5����b\�.��y	��;%�$I�P���D^�7N�����c�r�&<L(a���CR��E�H���!��Kܾe(ji�c��47���V�O���ɇcok�u��QH�l!�Ͷ���I�kV��q��yud�3}�}�S�u`�n_�қ-c��J�r5:Z���[���r�+�[a�N��QG�?����V8K�:Q�,ܻf n!���%e�˂nrCn�z;H1a��s�Ϲ�>N�?�gS	z��\�A���� ���\�`c�v���Ұ�ڒTN�q�Ǭc�SH4�}�Q�٭�κ�b�;��[��.����� �L.$4}\ߑJ�&��b��>�z��v�
&��i�.>}Q_��ΥdE-AG^�M�YT׶���Tsqڷ��T���a|��0o�/�<�������^�1N7��l���\-��@8�ߟ��w`ȣ"̥��g��u�up��?-�򝄥1����%�&��v�/�Dz/�C��B�4(���΄�W��S\��GW����呬0���Y�_��"b��F���$��BHmC=b�7���}U�=f�>?l�dg���Č�K��_
�RL����j@5�f�Mg��H5�!�j�T�E�3�1�Z�@��<�g�L￀�@Cv`<"�C�C�U�><�x*�4���K�<T\=�ӆB�ۆ%E�b�I�d맷�u�������>�3���Z;��z����2��}k��.�� =2��f��N/�"�'��7KR2@�d��j�՗����),I��K
��ew�Ru��������J[�}+�!6���jMV��7@SE]�9��~z���{$|��^U���@��ɉ�qHg�-22;�G%��`��c�V��>l�P\?_�W$�s��Q� �bƛ'X�&�le'��V����9�X��#C�S�==�3<כ2�v�SᎰ@�EWŘ}Ь:y��P�> ������"�@��O�V/�Gͽ��i��М	�>�/���]L�XaY��	Ł��/�ug0��G|��Zܨ��jH�Y����n&�U{&g��i�1g����"�aAb<�Y���VȖ{�r~d4�@��1o0�U�Pq�Ä�NR*a�u�J]^�E����G6KI�����m��;������ۺ5��۸T���f���6��B�:S�Of��_�z���R�Ɔ�m�'������	'�$M�����з��n�dI��KD;��Es���>f�[?
�AZ���'o����؃�S��*���K�G�}3�"��C-�U)a�E�#EU���m8�d��ئ%E$~��,���+{\a�6�^�%`��ߘ�o�֗W���M�<Z6��~�!@������a�Pni��AA�]��n�h�8W�*���GY�"͛s�z�wD��Գf�q}��Tܘ�P1|8� �t�R;u�W��ޯ4@��#�d�&~\��S���$V�l���	g�V/��ϒ.��%�P�u'�ب���q���<�0�Dh`'(�udl<SBM���R�ʅ��0������c�^��a��]s7B��C�~�6�O�{U'�P־&�`���Ʈ*ݠ�%Fw��n;JXAb�d����h����5����T��Jg�}�Uq�� ;�S���M���/��rgǀ����Uy������=)�ގ�J�f�+m�ǯ�ۉt~p�s6*�~�9�+��ԭݠ�qw7��Fc7�r7C{K�ZEb��7G��k��
6�P��-0��(�nM�|z X��ݲ�7|��L�T��r�km������m��b)Kj[��^�� S�,I8�5C1��zN�ǂ�mLq/p�6�|w��̅�xLĘ��2��%�hVyN+9��mV�l$�a��hbbl�7�&��Nfz��YhT!s��)V��W�������w���V8�E������Ř�L�h(�~^� �*R��:&����S�eY����`,~��j��Ur`��y1����2j�b���b�1]�iwe�eA�Lʜ�W�5:)T$[�>���E`���Ʀ������jN���z�$�K�"�.�h�l*�h�c<��<O��l���;r�eȫ�%Ǘ��H�_H�p6�^?^��<���[�gw?]$R���mcR2��w�o���ܑ2>��J5g߆i�f��pr����[4��5~*נ6�V�5�� � -#��v[��s����e�U@H^h>�=���0>�ʋ���-���C�*������=��$��$��k���;e�/D�8k&�����r��g *;�w��-3����X*ڬHA���;���W�	���`B�/x&ާp�BP������p`�?n�</:��Öa_��^������Қ�8[R]ū�l�̋����E�^O���>̼o�mp�v�]k{�=h�����2�&�7q� u��6�r�����7�o8�JO���ݥ���fI��"��޶��:�0o�z{R~�M_����e��l��&�+)voi=���f����qǐ�
.*@z�b#��^-�C[�5v��C�WtH��HuN�)�2P��� u�ܧOӜ� mt����\��qe����\��A���q��F�0��)��]�7�!����뻠�ѧI�k�>�⨌�3�%ɬ�,�rN��j1�2�b�c��])V0/��y2,�����	�\n���4|�r|S�x�@RC��qox*��@��!KUyY*�=B�z��&P��������l��)�.S��ۏ��m�k��7��51u�7!�z��(��Uz���D���o�X=*)��>ij��~�(�y7����]G�x�WMw0y�O�G���w��<�7p�^vm�56���x��� �nm��_׶�N����$��p���0�^�է����į:& �kϩ��]�E�a&��E����s��Y[z�vT�Ƿ	��������Ñ!Dp�ly�WY��C2��G���uX!�GF&���`���ڴ��V�x�����+�=��I�%2G���&"Z�(���8�ű;ڂf��W8�w����=CX�������������hW�ڊ��}�����AdHJ�M= z2��
��a�$�2�����x}s�����8�-V�wE����rr�K$Ds�^��	7<Ҧ���a���x@�;f�})���=�.���;
�����I:�Rm�En�e��s�J�gX�9�+Y6���o�f �(��K��uǏG/!V��|�U�7�l��8���*/�0r�h��`a5=�m�ݜα����Hr� �����\%��j�O_{q50�lf�A�q-��F~���Vni�[�5���-A%,��k�^����7A\����� d%���y� ���{��ɻæ��o5�olSںu�U����);�]��R]���:�����1���ń�	��VV��^m	MJ1�u�n�&�h	��v�g�#uכЕ�)4F�0��Bs�r\�QAp�h�\�ѥ�ƐґD�H&W(�E��\Ɍ���P`=���I�����5�;Ď�O�>�ЮQrѧ��&Uw#��;�(�[�g��0��K�������] �F�$�B���@	=vM�����lw�a�jK�(f����=�;W����b;ЁI?Q��n�S=�?�N�8+
�鈒}bfk�A�g��#�_�NS^�ٺw1A*W����
� ���}e @j6�Az���е���?"�2��r���>I�`����2�#�渚,�x�z����!��3uV=�;���b�! �c��P����k�'qj9	P��T僴Ƕ���d�Wui�l�/�
,*ƑM��M�Y��� -����E!i*�����&"�Ŷj�i�R9!���E��?i�5��us�\_�<��˿�E�1y�,xϥ��ہ���Mq��"��>��C�����n���o��
z$���p�|\vV��9���L�t�%T���b|�>�ͥ�!��>�V �U��7���f��<R�ǱN�Rj{�0�~�Ì6v ���6\OK���ٷ=j���9/���L�����GЎ��\�QK�.J~!.��6-�3Q�s	�l�6�eUܒ}R�yԩj����vԚ�3�γ�י"Ӳa�VU����� �X���~�U�E�F� ��z�l�!2"#�Z��NY���^��� sNQ����^�N/z(3�XU��U �l$0�n��3���|�����S��(��ׁ�R�&�g_7a��V���NM*�AQ�
����ܬ�l�?=�/Sj��|u'�(PWP�����QB2�R|�PB���K:�����0�]Z+��g����~�j#�[��������1��RK�(���ߌѾh��=/�0H�t��DߔܧŲm�>g�}��p���������-�@ֹ�(
C	�2�H�"ٷ��يo'}$��St܁�r�;����8+[��}�G1Ӏ��&�7��B1�Oi����&���P��u;�S��FYݔɹ7Q���,3Ʋ9^[��ޛؕ�ڱ"�p9
��m�of�~%��p�`���m��	��3�lOW]3ϣ+��i8�5h�ׯ�׫�lc��	���/�ԑ�_ڶ*j*�g56��r���NG�B�?���]e4��(�L��4���	���I�1D��C,(�@�ШN0��(��խ���w�f�P�-�$2j@���u���������A��eL���/�6�9l ��= �7�%إ\`P�v�[q+j=�f�^�c�j��IK�]X���ir�=R׏F�⬃�.�];�<�Ũ[�ɡ�l�$���7��(;n.f�32�+xK|�e�¥��� <tŨ�G~Ҵ�`cq۷͓dgr+�)eb f�%������7RsK���̀{�Q�'$,ˁ����W��d䢫T`�"��Nw竪ߋdd�Ss[��
��!�L@��SM4���/��F���wf�Ց�!�E��@O�o1Q7�I�
����f��.����;��e&�JIZ��or?����g���i�E��;$���yJV�z��ݍ����ey�o��SFsE�}����؇�%����[�K���T#B-�^7=�-ʦ���T�-��]�z�k��@͇f@�p����gv�1j�A�!j���L�W�?nM�TuJ�&)���r��8E��c�t����Di8_S����tA�\����K������+�d�
,����]�T�^��MQ-�>��`��3Z�]��9�@��b~+`j^D������7,L�}fe�P�t�� ��M��]$���t���;�&�4�ަ,���>����ꣻ�d��v8H�-b�"�m@'%�i��Eu;�P��Ɍ`vѐ���~&�L�n4H������5���f��𐂻ȢH)���E^�WK'��X/0��!�:碃�ED�7��TrR���(�{$0 5P��DT�.����U�P�o�6�)}�AZ~������(���́5����/���$-��y�Mʒ��*�q�U��!�7^όDЃ�9�"e�\���P�u�!�1����Q8��-�"�W�����"E�W�Wybp��N;�^�����T,3#�������ɐjX)Xj���N�8�'��(��[�%K�������;�>mpC� �q�}��T�fֲ�:jS�O����5K@���D���~����"����"���a#����Q�f���Z��+�������S6�-����<R�C���S$�Q+{n4dƟ\��{Ht���i+׮�w��$|Vc�V��E�[7d-D��.�lC�-��ױ���("(�ի�3F�S�������ž�?�N��6�>ޕ������'�{����	Bz�w��In79��.�(�	�Z�b7�.�38�?�LFY�" | .�c��|I��c���w"�����*"���dmȟ��qd���+����i4���3}ŤÐ��*����	3�;��)����9���c��nF�ֺ+�d��2i1T�Ϣ��;��w_��̒_��X�!�b	������q�嚁O���]z���߻6�U|9O�(��fa
ژ� �3K���>Άw��������K�t�b�I�b��C9G3�9����-����9*yY�����-�)B��WfcSO����3Ҏ��&�~�`�%�"7∭�I���)h�R|������ѫa���w-"ݢҙKm�E�jR�-�N����cT1�Q�ZZ��"�U�_&���z9�(��(O���T�Ɓ��7����c,�9s�K+�P��q�i�v���X�w�7�t��f/DG`:x��<m!:X��^Z\zڐb�hG�*`	P~�t�z]�?�@N��NALw�G���`��V@�H�	O`u�I��G�[��b��?���T 4�ZLV͹Gyø!�O����pT2���5ǂ5X���y���*>�g'�m��%s��M$��1�A�!�*#�#�7���-\U�ҋ��?��Z� %(�[��''�V�Z-��\^|�����>���>'��و�T�L���̶7��{ֶ�]���cm�����_�[*�t�K��t:
�4�o�4�?��N���b��e ,bu[�	w��V�MP��_���?;��J'8wmx��%���;�5���ƚ�
I�7ČF/b�UJVQ/wp\�I �PG���2��1L�Pg)��Κ���J\�%�9���~��(/ӊ(k)U�c	!p�`�cL�xݖq�N���!��3L=0�B�uq�~����Fe[��=V2�[�;��՟����z�_�u��7dE�6*ڜ	�+D�5�qY,1Ќa��)܉r�.�Y.�МK�ա/�Kg ��\)�vc	'z�{�m�����dJ&G~���DW�R�c 8�I}\ݙl��ixF�IUӾ�+p��Xtz܁oJ0Zϧ�D��P�)8(-��5���z�Lr�(�X �!�Icl%�����H��n|�eݻ0�%�ߏ<�]�a��-dZ�:����읕7p��'�좿f֧��=�黹�T�D>	�r)vqSW�B/=�G~�re�IU!g�V�O�+X�a,q��ry��s�@��yp���U��������[W��y	����勑���.�~�/#KTт?Փ~��������*P��9G�t	Q����}�R��b��`FM� 7��m9^�Q���P�c:�%&Z�x�Re2I�Vhzb��S<?�3gf��z��;F�oW���7c3�)_��>�>u�ײk��B����!r�ZF��s�P�ʱ�ߋ#������BU5�t4�3�+쭏�5!L5��r�f��ad���-�z
�Ǚ�Vvg
�N<�:��
f����L]�����-�i��<Ƴ��.��iv�8,�yk3I3�P]�7�'RZ%�\�2��n~�pF"��x���N���+��bmi{�ڙ�/�ئ��S>}�">x��}�"c�?�j^v�c����m[�����c�bb���v��L�� L��l���?\�HO/�Y��Y�Yq�`�C?3���ՈQ�چ����R� "X�l�JTj����X��>ų{��ʯ!�~�m�CL�0���>��w��se)���E0����m��[�CIg�K��_nC����F��Oޡa$ ��uO�w��-�È�ő`��Xf�J��"�}"
���F�ԧD��k�� �]�m�vk�d��$�\�]D�}� �l���F.DɎ[�����~����PX>p/�}M��I(F��-��M�=�[��2WQ���Dk�����x�;f��7�D����1�)V!"(�QA�3v�^�=���n������`���	��n%�%���k��7�Ā)�=?�~���~���>ٗ~i����o!R.��ǠY�Nn\T��w6��]#j���m\)�����\d?���$�;f�m�E�b�I��m�A�m�r�%�u�M��o�޺*
$v!����dԿuhx��w������c��<i�/�a�%����s���U���tG�3eqV���*Ï�:q�!�|:u��8%H��~��:m���ǂ�OIZ3�cT!����oE�T�2�3��.kB�l�M�`\T��_��O^p��/0����Q?��+���5�1����I�3�޺�[�~��`ލ��!���6�0¤�l�6#����+I/�-%�&�(_�!H'�����埰��[�&7	�`p\>?s�8�ĭ M9Q�i��,^c�,5�s���_/tA{UA�ؽ����o�؉_ZY�^X�u��%��X�m�9�^W��I�΁��v6����#H6�EqԜ�ĹQ�%3Z9Y����!�����|�;�@|d��(����u�c�p�z�1��6>Z)��H�uBw)��.i�+?�����@\�]sJ���M�qu�2���j�H�;
w3۶`c#�j����ƿ�~��Q�V�`�*&��%E��e�]�H�U�Pj�Ғ�ڃHg�dʱ�Gо��va��aݨ�MVQ�<�쑂Q�Pz��@a�Q]��xB�N*���]������-�1Ý��n�Lm��Ҿ3\oIé^�<"���x+W_.ِ���N�Lw`�3��=6;a.���5�XD��h2�1�@��1I鰙�B�dq�,xjnXNA���)Ep�~й[Y����E�\���f� 	���U+撏��;��_o�笳��cˈ�M���ׄ"��?�:�LS!߇�x�Π'�"�r@�X����3���9���ԛ��5�r�F�v���>;��`�\yG`\�:��f�_<#�l`Q�,_���"��T��Buo��aM�h���������n7+�=;#�YW1k([��p��
j�?Ϗ>{�a��B���O���I��.Kϵ��Q�{��T�.�{T����4/gR�����`�E4������7=Zel(W/$q
ʓjQ?�AB�Ud�-�9���#�m�q1�\<�ʸvÇj�1���MR�p0�hP��
Q�&I��@�23�:ko�C�1&��T�\b�ur��`����	�w35uo�7��v�Tc�����s#^���僻�����|Y/ʋZ��U��ҩ&����� �����g����,��Y���*�q	�4��`�ŇA�Kl|z��*H[uT��<�A(���XN]\�:m�m��`����T�5uue2�!��D����i<�ͤ��	b���<�R�Ԧ���ۤ@��}���M� ���MkMk$*�c�#���9����e�!4Į�P���\����m|}L����oz)��5yIi�xEYb���͘��n�A|�IZ��
Fk��ʋ<h��0ȫ�uߜ�:�2ơW��̸�Fv�V�fY�E�\
V�J}�lZ�����\�A�7�lS0��]ߑ�ۋ_RC��v��C���	���sи gp���*�)0���r�����Z��6a�o��5�1U^�]��u��aQvf,�M�7��	�e�e����*-Ybz҅X��k���Ѹ����䓦�\Z�R�v�m��єP�V �5��J���@�n]�A6q4 ������O��R:1�{��%�5�9 |bΊ�a=V��p�a�U�Ĭї�/r����b�*��t�:��/�2�K*X‬|��wp����'ʫׄe���O��=�Y{湃e���Y���1XV�b�yK~lue���\8-��>]]��W�<A���<@<s����~S>�7�|,}
�S�Q�e�b�sd������a�-�hh��ig�,�Q2���;
O�������%�D�<Z�`p	��z��tΙ��"u��Z�O�ʶPR�w������`<I���Ѥ�6�Z������3�!*b9p�`],o}rRs�p�S��l�l3q�;�|4���_!��$&��pL����4d,������R�`8ii���>�����1?g���c����:[�z�)
�J�i��Z�$$7Et9���l�8���}��z�@�Eh��͠����6l�{���PY1�Ց~��Za���0�F�l]��"n�D�(Ťn7h��{�v)����UB���)Iq5���V���s鱿���AD��e!f�xƔ�p'��T%u5M�ہ�� &�ӽ�F����A�f�7>��4�����F�ɓ�O��Q�\=�\Փ��+���m"����^.Z|g޼TGn�����S���p	B��*��l�V���>�Y�~�=�,�n��N�m0�A�j@��|����Βw(
��E,s�WmuJ�9/�W}4���@sc���R�_V�?XM��/괿�T*b���~�T�:�0���Z�Kz�� �=�U7у�a�i,�t��v�XPA��'��b'4'��4S   g�����r!��۹�cϯH���>N"���^��h�LU��q���ȁ1�gI�: ;���u����/�4OC�g�k0�հ��NX��G`��n�k6���X�hhdocF��/e�![U�7*g��183�ȋ��)L�l�>��cz݁����p+��Œ��d*o@��U$������L��2/�V��( Pf)�<d�W��wZ�:Y���4$qed1���������/z��q�*��W�w-m�/3��R?���h!K/��˽���-�խ��J�P̎)���0�ZJ��ri��'{�R霣�bčUq�$[�>ud�/�ٷ��΂KH� �0t���4+W^J���5��#�gi�JXyP}_�������C��F��ҏ��ө'b;@o���{jB%G_���;ú�f�o!@���*-W2�������&DJ�ڰz���]J/��'ڮ�{�!P��P�"�d\Õ�\a�~,��V�%Fd��w��W]����m��l�0e�0T�XJBk��=��ȼ�֥{k��1zC����μ���	{�
x��q���s��(P���R���NB�M��)xe��$�0��>, ���aN��]�fҍ�G��0s�'/�F1��iH!�.~�`#��0���i���-ˌy��3r�����f+�9U����̾l�|��?��^�w�{���9-�����ln�d[��&��g�uš��]EC$��C�˴
(\<Lyy~�����W�B���C�^�^л��!��������\^��'GX�9X��SlI/�7��L�Lġǝ��0-_�Ńz�X�3������55�.;�t�mYh^��5a�4C��(��ؖ��3�����R�����w��JQ��=	�#m����4�� N v^F5�Е�pS�x4�����$�ß��:*���DFq�{��Xжvk7/����m�|�����X?R�((+?}J���Zֆ���<���6����M��.T`m�PWF8��0���N�V��kaJϏ�$��f�@��d�ē���OV��Qo��d� ����se����C�k�yHR>�e��e�V	�>�~�szYj�ȤΧ͔Q�'�1�^�'�;�N4�Ex��[�{t�EL����:�N���Ch�3
.��Vc�! �
�Cqɉyk�-"�n�X�wE�#��p��]�gGܔ�:�,�L%���2orb�`&�^�����47U7N�ȗ'�y��Q�9�J�w][@m�n.X0�������y���p�=A���×N��
��Ѽ{���^�zʏF��7�������	0�p�̈�;h.�Ӊ�5��5K�)K.=�/o�`�E;�[��i�|֛
D��]��=*��2o�jnb_�2h��n�~�/v��}td�U�+��r̖2&���J�;{&pjQ�@\���I{(�(��!�o���/�sǳ#���oM�L���a�7c�;�"���E�v���R�1ƗIdf�V�4`��H�KV��tv�i��ځ�ҫ(����.T�5�7�!���{�q�1(s�&]H�'"C�4ïB�E�����W�z�A���9V�}_K��?HO��eZӅ�yH;�� �QS�$IO�Q�֜v�zCSl+��#���Vu��AΓ�#��|�X�2'��a)I�U7/���L<�r9�q��cS����_�q��_deӣP���^�"p�@ar�,����ѧ<� 2%C&x�4?�k��ԯ��td�2Egm�  o��=B�N7�)[����FKL�9���d/xxd�uѱ�=h�޼,�~1ď�߷a7m@a��_�e�bxE��=��e1��U��ګ�6����Z�yҹ�(&:}�{��H��b4�����<M�K/�nZ8�y߷~N��#͋ xØmaoke>+͞����7����x�g>B�N�2:�$<m��O�_
��R��rVTth��ݖ��ޔ��"}Й:Bҋ�3�^&b�[�������?���*?���3J�s@�|�w��kY�B����U�>M2�H�_m�kOD���Pc�O��2ݴt���u� wS�$���w�3K���i��Q5�(k�	��tP^d�t>P�BS��K8s�C�����\������1#�� B���D��b��+WP�MZ
�l�馊�ӯ�S g��uʨ�?<��Z��
N��gezҬ�K�$�sD�Us�s+БT��	b� �N$�#׆��o��-JOwn��7��Ѱ�eg����K��w�Xv�f_�Eꝫ�� �Q��]��&��B��o0������YR9J�N�n����b�<U����G�[]9;�[}�Ų�z(l}���/���!�E���u�c�{���:�0F��ft�zBT���X�6cYǴqy�I.���s���=g8(�m��SB���A�z�݄���#���/>���C��س�W��Ra�o���]�@u�-`wK��ī��7-Ɂ�U�HdL��Luj�#:N�WBE����f�A�b�8ޢm�O�%]QL����&�����;�C>Đ�w:ԞU0L�����i�MϲG�t�ZsX���D��шK�-�ȼ$����!iI\v>�n8�zK�b��T�.&|�i)N4,柈�w�������FJ�0�	���%�Ҿ��SZ� W|�>1D*IKF��$�u��(ɰ�x鋤#52�a�k�P嚣��M������ۋW��}=O1���?�R����;�w�v�6A��L���_�N���؉�G^��ۨf�-�z+SG�Wt�%Qvr���\2O(�'�yW7�m��u��Q�9���C6Ww��5J!�����7���?B�w�~�Q�ru�d��?������N�>":�gD.���,.�F�3����_5~6���Z[&�"'&�j}I�C�[q�im�C��É����_�y%����-恔�N���D�g�9:P��F����T;F�kc��8��}��`M)*���Ǿ�Z�$�����Ɵ�S.�(��߰(^:�w�?��%^�d��ߖ�?w�b��ι�`��ʲ���s�SX��w4�7'r@��/����|*mǩK(�A�\q�i�ߘ��>>��+h�PdQ�4���R�Qo�R64X�&
��=b���i�`�{s�uJ���=(�~j�D3SK$Z�u�,m0�Ӥg+"/)�U�N�����^r^��]�Lnܵ����Oܢ�N7���3-�e��#��qy��n��<e���P�:���"��6����jr,{���*�u�[��щ�K�.Cԡ�ٲ�L�E01�
�0�ע���; z���/�����/�3q��t������d�S¡ɣw�pO��/����K���# ID�<�'��b_<��o|��R@�tv �rl���b�(#^��Q�2>�/��ʘ�9~x츹�C[�\�銆~>�W=?���1���X��bO�U�^�1�/E���ڼ5��^*��O�0�^x/6��8�.o�>�����ϱ��w�����o�f09���v9��B�>E�;�����?��<�킏�jD��e���;F`��jVxC�՞�沤�^cO|�����8���4.P]�~��V�]a����n�����$h4 bX}%��A����D�b�M=�?I#�g�j�Q���]�ө���::��:���k��$�M7ɼ��ԜiV+1a֮��gG��F��cT6Ys���[# �,6�m8��=@��l����[`�(,"$^������P~���YH�J�S����{�h��f���<S�ϒ�%��8qsCl�6 ����s��g¹�:��&g�si�J���g�/5k�!O=�o%��(+�.��ê\ؑ��S��2�������� �q��@16����ml�b��k�'a3ϟ�#��h��d����=�����ʵA$|af�$�S[j�������Š����z׷�����Y�O�]t�����inn�d��ZE����yD~
%rr�a���S�Ba�]u��
\S��"�2p=��@�9?̧Xރni�W����ğ�2zj��b,�Q�G��!��O^�t�N�9��?J�o�@�(�N�7Mٴg�>���(�6��kz�GV�������}�TW��oyd��6�p��P0NA�zH�"���(�}dˀ�LA�O���	GغyÉ��6s�sp���(��՞J�R˥초����M���#�%��+��Nr�MGՕK���#������'��	y��Qu�3=�m��"X���l�5�#C+/�e}�|�7̿WY�ˬ~q���OCH� �l����v������^��籝8%{wPM�&1@lԫ]A�i�4��t���罴�8�On&ߘ��	m9�Z*����Qp�`�f� �*���TT\��8�FL�� ��$ $�7K$BL�=F�-v�~�v�D�'�^(њ�O�H�~p/*���.[��SJs�@���ü��`!�|ˢ��e�pF��:Va3fʒ3O	���tmt��̀*"���=d�~�j�[�����y�5y�2�6�--a�6����D��J�*�)`-�!���Ƀ��U&�S��EԵ�JI��W��u�x���j�:���aBO	���q������c�;�Ǫ��غ��>��/�X���Z�CF�h;~� q�!�I����9�%JX�>�nm�~q�����:24N�����Uu_�B�����,+]�3�=�ż6(D&�p2��s�l�D�A�i�H)��'�7��5��u�k�������}��'�*��.=��h|b4gV
A,�د�5JP���
.�!��	GMK���W����E�tGӂ�%x�pر�&�� ��B43��2�����W�}�
;�U�7�pM�������f�������T��rQs�W#ǘ�r"���(Ǳ,}v��Y���d�<� �l]�}$��j���t��@h@-,ޥ��u��]�W��g@��r��_�zou��Y��*G��ͣ�3���uˉ$띖!�gf�L�3z�v;-F�XW�]&���IE���c�"�������_7��N����@�-��ׂ���}�gݜJ	5 ZNi�}�k�%6W,�'+�H:��'X�z�E,0X}N�Y�?Ss����u��[�C���@n���.��{�Bβ2j�ҝ��X��b첵l�F}�U����kk-5�Q��EeY3�^�_<XA�k��>6?,������ �\4��M��+5����[0o����c*tw��h	do-rq(����o���H�t������*J@/�0���5�I����%�E|���\x�\W
7'�/���8{�D,�B@j���:����Տ."�ֱ^ �(��ٵI:ˬE(�?�~"��Y\�eQ�=����P��B�L�
�%P��D�n������1��7��g�?�,�L���0i=;���U�o���	Q�b������?IA�Hr�m�y<z2�,�K���dB%���5Ml'_����1ƠV�.��jF�DFD`�J��*/EUʄ��͊���XT.������Z�j<#�;�_"�NG1�#~:}��G�9��v��I���@�Ϝ���e�T�s�o��B��mu�WIP���ں�^>܄#���ʿX�Ř�.C	��Xf�8���?FVr&��᭍��
�^�U���݀?s�/�L�S ]����t��ՈRA�g'��>� 6:�A`����Fs�f�_����H�|�7O=Za��H��n��&T�⼨�	=���[�����*�;h\�qZ�eyV�MB=���3�����,eNǣ��dM�|��ui�"Hz���w�ڭ)gY*_��Y*fiZ"���H����y[NL ��h}nn�O*�x�)XV7��TP=�,��o|���<+F���京�p+Ѥ0U�THJ~G\�9�����86��8Z�C�ȫ�"-���P�R�����3�����i]�`ޞ%�S\wv5� V��W2��!��[5d�U�)����0"b_|��lXJߦG>R��(���q]����^��N	�X�a�[�e�>)|Xy0��*��d��=�&�L���&��<:i�ɨ���=ec����0��!�%{"״���$���������5=����c�s���@�a�/ܣ��O�ɬ���e���^�L}�A����X�mg�M$%D�<�l�D$�u�/��Ӆ�J�ܶ�(
����3���ض+y�+�0�tG�C/ٖ�+�� oƎ�P,�*ba
*]x4����u��$=i��y1���*J�����{
���C�\r �ݽ	~��܈��Ш�	섰	9Oi���߸nhfX�ȩrG=�'�s�<���d(�!F����S��}�@5���د��/:�~d>��B�E��N���9�ޒ%i���;��,���Lx��R����yT�en/�A(�v�B� �A� �C\�S��9��A��3�����?*>�9D���T���A��\Ҡ��������1�J��,v��h��c�8��z���5�;��-��X�1�T��o���Y��I��Z����ƧЄ~��q�b<+4'/;���nm1����|6��?���Nێ����=�hV�Z���c�a}��SI��L�U?$��j��йr�������R	�ǭ�]�e�6���CM4#�F-\���VvfD�����q?fJ�hf5"�mp�
��-�lf��z��,j���X۟��D�v��߲Q��g���K���@ݩ�z^�/k�/&k��TZ��1D�n���W}|���c!S��D���zʣK��,�Rh�_I��#ؤ���f��6�K'��v��h8� V�a�H�I�6P�(��RHvaYow�����e ��_'OĒ}$��I^p���q-f��7}!<��J����!�(۵��"��1}��}��է�_��7���[)��L�7���1�m׹|����?������٘�,��PĘ4b�d��Μ�������	aI��,]ۙ���2 �9�g)ٰ m��[��f�߁���z!��:���~o�qwz? 9�Je΃��]�4�gn�t���m~VAm�?���M��\8F�Ȃ��XzL+d�K��dc����$킙w�8����8��A|!�k��+�a����b��T��R`jZ�#�EM�����\��=�EA��C�D��1�ݩ!��=
��a�����iw{�­P������^�qb+;d�,��2�{�*Ag�S��A���@�!���<��q���^T;ƣ�־6D��cTq?�iǤ��@2�[fL˓9�u�w��߲��!҇�_�tI�v���H��v�Bߣ������/'#&7����Q%+��O�w��0@�K-k(����g���u�|�y�.�Q����G�����.�s�D�{;��!��u8攛vL�n)���YWug��4雎�\V�'��k��[��t��
�W�m>#5�6zt�)����q�{"��mj5�6�"�^,1��͗�b�_[3{AV�Mp2z�J;$?<��<�
4��g���_�y�<�i�V���Y�W�j��7ND~�=�M��Ϙ�X�
�I��$I�Ik�����{�����J�b>�>q1����~<���;W���a�F˷��ix�^	O�S&E8�Z"ۼɡ,�g�:�L�Bw�	��p���D�~SIN`E�ޠ(���5�{H�����FL�Ӷ��#�&眤�g���������_y�Ħo���;:���%�K#<�����\���z�癭���Թ+�yh�acv�vk������&���܏��VS�m��8:;6�_{{$�g�u��x�
.�w��ӆ@y#���������Rj44u�iZ����&������K��q��x	�1�u2�]R���"Vmq2^�Xl�<���=~qQ�z�� U	9������*E�X�9�c�m�p*�gSFj����h�Ϋ+J*��1^�~eGK���ؙ='��)3�|�/����3�K*�8�1��q]�����.�~�g�����wg��]6bY�����W9+���֪m��L]���C�V�tS�o�u�3�A:gm!��^�M\�]��:a�qj�O�I��&B�%��DTo� ��6
���gM��i;��[��a�nYt3��9_�a3�(A󓘣����М+?��f]�S��8e��ϡ�+�s����if����hFlBݜ̶oն�������|��"�e%�؁�޶��l1��S��s�Aʋ��W5��>�ޚ\M:�V�C�.g�:PR���_"��·��7Yt�"#��/���� h�8���q��i)��a|�# w=��W�<76�Eng;Sڰ�M����l�b��
�	�.�M"_q����m���)њ5�����zԌɯ*r�5ne��T9��M�����6�ߌ\Jr_Lxȕ�D}W�<�������AEԲd�����S}�P�\�"�Yr~���@�Ĉ���R���I�XI��+�y�!�D0��u��|��3e�9�OF�l��w�j�Yk�T;�h� �s�
����ܯi���_ �1ʏ�ڕ�=��� �3xF������~�6��v�b�����J9ۼZ������CS��6��Yh��󦹹��7}��ؓ�5Jԭ�Q���|�x����A/��O��'��]�
��R=f����^ȁ��V���V�`>��"˄,6{��
��5\��I�H��u`�:�E�P1'~#fe�-��й4d��Tx�+'N�
��ƆH���Cv����Ȝ0��ܷP��o�f��]}
�7� ���g�C񐛫���t�'�r�o�ߵ+$k��ܕ�}4�u���ҍZȞ#L�N.����m�|72٦����b��8D��&T��Z��J��h��SP�Q;KX�8��r����mB��g�YJ�2������X֤��VA>�#���ø!ȯ��۽�+������m�&`۸�9u;�����蟺B侧b��6�"��m��%�c��q{b��mE�޶i^��B���&G�g�L[����8f�R��:���W�Bf���v�֎�zֽ��AL�{��c�ԝvU�>������N.��.(�6}A!e>���q�V9p��wJK�+e%޺l�h8�弽MY{7)�v���VN���&+�h�|V-qx��*�$yͦ�V7��!�l��X��)�ye��T�0�5��T?u�yi�4h9��$[���H�Y+=<+��=�kFR�,�T�����9�׎R�x��r>���@���y��?���r�S��&�5*��!*>%�]y4�G�d"��A��ǷF�*����ݏ@�kK�i�{�*�j���jce��h���a��B+�|�$���1!�Y��"���
��<Fl���S�ST�����'5cJ��V�մj�4�dHC�7�0�yo�N��X'8�Ɲ<߃c� FH��s��ߐ]�~�$^6��>�(R4��Q�߻�G�1���^��e�"З��Mxq@�*y�ߊ����=>���̨�i>"�s����BH�°��9�o"Z0��*?KqO������GfV][ZzU�M��'64��*Y�f�; ɋ�޵��C#v�p���5�7{`��;��̄�Ս'\�)pS�������7��a�g�P��"!i��+i.����!P`����]�_ָ�z�#��X��F����?�P�u*m��;I�p��V#� ��*ԋ��_�3sn�U�ɓ���\&	o�1�oG����&Yi{ԇ,�:�I����]���ܴ��Tc��_��QMg�1� �1��z�Av����P�v`�Lr5Hk��'Z�	}�#yx��ɬ�s�����=��"%s�T�U0d�MF&C�Atɋ:����A���fE��w��6�}xv��8����O�F�>�<T/Yę�O��ieR;����=4��I/��DhX�>�ڠ�B'�z�cj(��2ύ��vr������'���`�$v�۽.0:4@u���z����X�f�a\.w�_���b�%�|���-;%/\\�BC�>�7���.a٨��������T	��58ЙYc'������(��#E�`�ծ:�*�y���=~�T�.��Y�HdG@����ܺY��<˧��g�<y�̸
�����\�ŀ!Q��z�4��&5�u�������^���w��9�X��`&/�&��Z��ٗPx�[�)�\�
5�C���]q����-9�z�vD�2a檙 ƕ.�"'0LP_�����h���\��_=���b�#�~;�c�X����=A�F���1�������s�3�M�f��5��B�A��`^�Z���k�iI�R6	��t��6FK���J��f����ݱ���}?ݴ�s3�J-��{h�Ԥ�rW�	3Q��l-�`�6_Ɓ��m���%�ŤӚ��p�rlg�M��W�C#n���a�Z7�h��t%���+��YI��m��LbIʚ�=��ѫ�^@!��������Ef� �65W֩4f?*�1݋�x��R$JƠ5�T=�ea�D�Q^�R�@-�����H�]�1�9/�|9;J�cM��Ī �|shw4�u1��x=g �ё��{��d�͆�2V ��֩��'?� -fzm�N�0b��n����8C7�C��>#/@�I�*�?�f�8��1G-�}Z���l�yzaMԓ8(07���B�oC^�f���P�������d�]�|��a�܃jswx����@�k�o�u�o�Dl��B��Ʉi��}��E��w�@?Y�������3B�\6Pw#Tڟ�#R��/�m���4=�%�fe6�+	����Ӣ�ܓ��ҍ����$EqL��i�E����&$��@���i�����nU'�@��*jL��i`	�� ��8oE��W��=��=ln�drڇR��36����?�m�_�V	�"RB9h��IQ�znòy�y�F��J�o̦���w���5k�4O8tx"��~F��+��	'��@�����7�j�c�،:"ã�#��g'�p[#jЭ}B�@x[��8�f��_$Ή�-}�!k���d���0����kW=!t$>E�WVM�UIڧ�
��6�f�kJ߈�4�21Tײj��=榜�d����7��g��QN�A{�Ul1o����
f4��փ�l�,n@���Q)HF/�}�.�z��	�r�~{H��Ĳ)�6˲���~�� IC9����t
��O
#��(ɒ5+�p77-�Se� `<;���������[Mv<B%��޾ ����b����e�.��
[�X�q;�$;�1#C#�d��AR6
��Hl�j3��nQ`�G��2���.���D��6m��q�"1	�3�X��3�3e�qg��D�g�`�zs��猍�ա/���!�:h:"�U[8)D$��N�GD�Z�{�����Ϫe[���sxO�6��b��f�K�fl+�%�!�##��8:�1�̃�V�<4�yVZk�S���n����!�a`c���� �y�Pzdm� Y�4�;]W��0	��5�1m> �+Qո*I�a&�#b��ѹ(�ꈦ�k��(!��e�>!��{;��ptI[��#BO=X�<v����}����u~[����s��_}ٽ��J��9�t��[��ǜ���"=�D�V�(�W��s$�54q��&�fz�,IQ戸��4����ؘ�����F�p�]���N�5J]稀]�+��`�D����q��3g���Anr��7���w�'+�XU�CqZ^b�V}��}�%�Ҫ$"M���!�i1�Y>�b�\�]�>�jԏ�Y'���IG�R==ҵkq�d�E�I\	w>*W��x�K�cje 4s�G���b���/�m�u�SW�gl$\�W�Ȭ�|�%i�Z�v���S|��VL$ u�To�$Y��
��{�ӣv��Y��lQx�u�X��>~��n*�M��]t���x�n�73(`V�`������+�9��b�����a�P�%Mu4�6�Ft����U�v�7y�~��1gA3�m��ɯJ����zݴ
ܕu2��gs�sټw@�,6�\-U��v5�GZ���OjH�7$~5����P-��I��d��d�N��և���Ɠk����s���b�A�p�o��X�U|s"�s��H��sq�O�_7�T�̠�)�
��7��I����b�h0D�Bó��_�}���:p�x��N؋��PB��ٮ���a�f(6��YjWL4z;_�T�5"��gw_vit�T�ໟ+�]�Ub�D��zj���I�p�>�%��ɀ|�/|0��x��߮��lP��f��R�(��q/��`�)k�x�O.\/kG��W'$f<����>HV��c������s�:��M�IJ�ڗ���x���
b<�x8]�c=t�G�A�
9��4�����RJl����4�]�μj��͒h�J����ब�DV���`I����rCH䀳���0�5��e0�z�Ӫ�k�J����/*�ި�&)�h �n���.�ۉv��rco��	�QA/±�l�� ��۔�{L_$�O��?'��v�"(�f7�9k�C�i�C"(��`��PMI�%�|b��3{��[���%E3�_@�Ux5�E"�?���ݾ��EB]8�� ݱ�!�E�xdS�6�0�(�e�x��A�l@�6{F�Ë�A�y����}����7W|Vp>` �A�m���:ݕ��C`�2m��7�ų�=�R����}r9l���1�C�D��������bF��P�O���.=��j�t�MqF�_$�!�j\iaiP㢾�mO�[%�~6���y
�J�01�[�#�b&��p1��վ�9�\� �K�_�3�\��$���/5�-	�0I5���V,q���F��LW�SC���h�.Y>a4�z��P;��Vl�6�/F+m9S\���X{�����X��X���U���^�5�LN�AX�v�2g�8L?��aTMa9S��]j�.�;�% ���q1�s'=jw�Ѯ��禅�û�,��o{�I��%r�� t��r�`am����ѧzDx��P���+@���[,�E��=Gly���h�5~hN�[7����� ��]�W�q��k$�Ejo�����dC�_�B�f6�$@;�C<$0uQ%r��˜�xz�k����T�=�u:g]뎉���;f��-�6���v]/Tx�qJ�НH%O��D��dB-ʧ��ߊw�9�n�Z8 �Vۼ@ˋٱ>�~��e�wY���P�Ư|U}�C$���
�y��F !����A�GƠ��4��`.�*5K��qV%L��L�ܼ�p�b��l��K�D��οUZ D� ������������[	R�ʥ�Ĕ�^���՟�d&��/61
�+�g��t�y��/���)��e���ɟ�b���i�dJ�@^�֮D ���G~O)	�S,�:���wH����G�	�)���Y�<���T���S��o$� l��
�Bx��A-J�t���i�n1���ǐr2xn�Z�f��$:o���Ey�_���
�|���D����Y�'b��E^+HS���h��f��k�;��ix��i�S�i�x��4�8R>�����8�^�0�����^�&��e�'��-FL�Шg�K|��p8\���G@bDΪ-ۓH����`Wx���P)���l`}�8p|Q�m�P	�&c^9�%y�����_���h�A�$;��F�Og�����ɔ�i{��FjkM�}IG!��t���ײ�����X�]��P3�X��RD/f�G�@��[N&�C"}C��-��>���r=�������.7j�F�q�<��/jM�	U�j��&����F��uřq�'t�-��-�=X1�X��vdo�_76Z�c�]�ʉ#{x��s��:��tk�rd�4Cy�6�6�uL��zPON�^���[72�$���٥2��|u^�n~I����Av�v,Z��ݖ��Ch��A�y��$�� .��R�pɗ��@��U_j$��op䨇�c9-2��k���R�����rb�$��/��� ��B~ر�%�&�l�['D�c��k�Y�v��F)���*H$���.���C>C6�lPi������	(�D�$j� �&�����9�5;r<�U	�q0L���p�Z<�V�K8�M7�:�>b�k���;"v��ȧ�ԋ��	�yUI�3��^�-���<����"j �U��Th�#���MXS�IQ���Tb�~��_���޲Q<�!IL��L���:O��#�>�M2��嘺!h!��� U�+^(Il%�K�e�fe���ce��@�)`�Z�g'�>�^}c�1M�M\`�tER��Kf�A���@xڥk�	�9�ȭO-3g~�r�;ۮt��(�|�E��¶>�g�Z}(��z.�b����Z�Vz��3���ЭSN���j�l�}�5�jX����ky�6���J%0��I�I{4�H�}��0���y}��%�]�P7/N~Z�M)��v"�:�f� �t�$@ ����_B�̚K��a4"�����C���W�I���32^aU5���~x�9JgC���H����ٮNǃk0zR����a1��ا�]��oZt)�����f�O������k:+�ڄ��yq����6~�&cZ�u�?�Ӭ\@���|x[#��a��� ����b�zD��B�S��?��1�(1�27����Tz޸%�^y_���K��[M�:��y����`�cF�ܑ@=�,3DQ��b���-�oF� �%u;�׿����\>�y�O[���������L��Ako���<^{������>L�s�����ԩG��k��m�z�=��5A �5���aI߻�e6�4��S�B;�۶DdD򡚦o�[�n�u�N�x!(wU��=�����E�n��﷥6k��#F�$%�E?��0��ʝ�i}m��8���:ˢ����1ϥa�����J�KJ�Ú�MVE�SPU�o��}�u>�E"5@+�|ժ�_4�K��ޫ�C�d� �
 q�� 4Z:@˗r�_2}����N�{rw��&�R�]UV���<ƭqK5��'���q>�W$�6��`�˗�t�zc�p@t7�+���G��4q��ڳ��2�A�}��D+�cןV�Y�|)��x!�i�<ݤ�F�#E1�\2�ц���sV���HAT/�4�Y�Fj���s�d���-T�F[��-�^7�x�C1n�������g'�U�!�%�A���)�����8rLdԵ�<v��y���Ȝ�>c@��G͓7[���a�t����;veu�&L�]�q�*<?*W:P4N�W.�Zeu��l�,�h����r'�&3h��������ii�|��G�Ơ����wk���S�Ơ$��M��o��{NT��dpN�sJ���c��
�3j�k�A2�N,-��o���z���2P��^���`bB���������<�]ObG9a���F e l!�؅|��F���8�oK�w���a�珂G�K ���؀��9�m�2 ���z��J�ed��t`%�א}��N軸So+4@�ʕzN�����q������k=���;�����p���{��ۧ��:�z��G*�_e�Y���f�B����>�����&�T�ۃ�^��h�@پl�<Gk\3sI=���{s���g����NL ��f��-�C�G��rP�������yWX�$����l�DA{E^��
����{�n�;"��6~(Uܻ�������y难����6ɳ��U���5�D��KA�)��po�}I��|�VuͿJ�s���B$����ILk��H��$L��m��R�����Mѷ���NK֍2-6�~����>9F��E�tǧF,�HBoq�r��/�y�'��q�����8D�� �6�>��cAi�P-W<W\mVפ�;J�$'㟷�A�=b`����C$��t�Zu��z��R91�!��"5Sg5(a!2u���e��u1c2�ɱ�|+����c�]
�3�W��"D����,�����!�P��#5L+<o�ׇ!]��#t��J�,�4˝[2�P��#<A�A�q��D �}�m4���~������W�����ʞa�0�0�W'���[->¤��2��v�Cr��.�ō��ݚF�l�"Ԧ��e �@��A�
�MF���D�ʣ`�'��|e�m��})ē)'6V��r呯�d#kXbN�uB$�y5���5�<x;���	�졨Q�[�*���v܈;ժ]�6q��o�����Ҩ;�琉��3ߤA�� ����tp�L.��\�[�L�V �`�%�!,R�)�뮉��@��ɽ�{������!�{w��w��f��V�[~Я��$�\f���N�<���\����~4QX�B�.,��l�j��?�� ��-)X�alwբ�P��E�w�E"poI�c�S�no?߇��o���v�`V��zG<��[fElz;77��g�Si�Z9���t�c�5N�_Fy�>��b���Y�v�z�
L�Ѹ��� �6z��::�=>`���w%�5�T�3�1�+��lz���"�W���l��:�5	��? ے�Ó�>?(�J
7UEe%��9RE�M	z��^ �����E��$o,��/h��s�R���-��ՠ�O]i�g��.��m�D/�Zo/���ͣ�'܌���l ��q.��K�l�W�2�qt�0�El���nk%��Pm7��b��d��s�/�!�"��V^���"���nP��I�D���N�Uh�wn�.����Q�8H��9���2�)�Wmw��������7 $~ޣ㚦��l��z�q��3��9T�iB�SR���G�ѕ|�}+�ծ�41A�I���D��(�륢"\2�5tZ���Y@��<J͟J��K�l�b�J쳣b�i�����Z��#�ҍG೯=�d�w"�\^��PN+�K���ή>rɝx�[����#޷L��\�F���w_���+b&b����=��g?�D�7��-��d9獺d�;z	��.k�P�.d��e>����;8���@�C��W�,��%&wWD��p>�mu�G�1:#��d�0��8�.��X���ɒ^�>��c���-j;߳K�ף���dp#uwو�c�� ��c���}%H��$b���$h�A���k�b��0����%^�ǀ�)����Pbd�Dɒ4�²�1�]������jν��Z�@��w>�QͻexJkM3:�	0n���1Z�M��,�<��X^�5�zY�c� m=��B�����T�r
3�1N&NNd��[�ӷ���C�-�w�8��k��^^����&E���X�8�-c���ؘlZ�@ 4O?�d���Z�� +���ױ�]�@Ğl��JG�"�VEV�."F�G&�i�r�^�S���x��q�S�P<ɽ?�2��>`�}�i��fe\�{��	���î�Z2e9��9rdҩܩ��D��)��+�cmHJ&� �H��-�y�c �UN��SW�aQ�^c�q�90;(X|ͧ!����g�Ep�`������I�!��- t�_z�ΐ��ɕĊ���������N}9ZY)�������ݙ6����͝-��P��o$��$��6y��i�����}hC�Ԡ�r�4�u
�<�m�t´&&l����:)�_ԋ�\���\,�|�����I�.��`ړ�4f�i�����ծkHČ�ā��/xX0����>g�Ug>�J��ܐo�R��no��g�vV6:e�%W� g���Q܂-�87}�?����q@��VNȈ��F�A3��qXx�*ꊅD�}+D[AcO�K���s+;I6��̏��O�����˼Ϸߡ���|9VO����}[�[3{�=�ђ��dx�;�\m��]A�.��J��:<���A�t�w��AMC�CH���;y��[c����|x��XZ�'
�4 "�XO^��z}�?B�4܎�ī*����兇"��І�T ��+��]�Y�O���pҴ��'�~R����d���|��fA>����M��ba�G���"��dM�߇<{�
�lz�p���i&�_�i�oj-Y�^�1n��=������H�+˯Z>T���'u����,G�}�S��m���Az\*�jV�s�K�5px�����+6�Ž��oҡ2���f�~��R�2�2���Ԅp�-W!��sϾ�o��h`ǼJ��Z=�w��#�X%�1/�en~z�%�jP��iT���?������M�T|���ʫB.�;"��ѣ�[�2�-�޼���f�Wy1K�u�����^���,dbs���Ê��AT���F�9N�|���$^*ou8Y��P�X��׸�	
�f����zpb�H�;Bq����ް�*�����l��/*��Hi׽���C K�Lr�O�R<m�R�܃ɓ[��Ro��� �wB�]e�0�)L����A�4UbI��6\J���&��MTxM�]EN=A�H{��F���͓]�N�*^���X�;����Nب����)��6l�ȼ�<�nr��w>��1�`<��˦L�m�/�9:i����V��I�#6؛��r��HNX��Hαښ8�����B-|��x�`��E�$�J" M����3�'����J�8>���׭C���ѣ�h`E
9 J<��w�&^�w���%m��QE)����Ԓ�ilgR=�0�b���`�J�=L��u������ə_|�H���6������EA��2<&�Zk.��T�Ⰹ��\k,�N'���7���gd9�zVkEѬ���u�0*�k�_A���u�������a�mDk��T{ʷ��'J���oDc���3��H�>�%QQ��3}�$!�C%��e���'��nb�Ai0�`_F�[<R:�iC����1␠"T��������e%�'z}���2#A��8�L�̐/jY�aD�� ��(n尲���@�Q,�52S�x��7a-�rSW׳l0hC<�F���i@�=�������[U-w[� S]�f��zQ���dZA��ZeF�_h����p]o�:(f�F���9_�0��d��b㭍�3]&L�Q�.>!����Y�pT�'���x�"�I�cj���#)��A-�8��|����:>	B��ᥤiQ�km���E-<$�w�66��a,�P��!7!2��#��ɅwU���~5��w�v��/�>'g��=i��?K�}Wa��I�v�S6��A�<�ݕ�����x"K;�,���֢�0 �YH�%8��UruYVz���Ч�%��y���Z��2��2Y�%lcN���t���VR�D3���������T�h�u]�?#�[�p��������-oK^�j�ᜪ�K$�O䉬����^���F5�,��@�U�C��NI�ǧE)�F��^&���򂒧����w�n�f?-sǷ}�{�t������9��8�;���C�b��nt���-��싶��fF�-�'�U��9�$�(�X܊�sfP�:i���Z��������1�k���C���ǁ[����B��{�6�)ʲɍ���5=�P/�leǧ<e���0,�g�
�q�U?\E�
,��	�1�������aI�M�<��$��npL@O2���6GF��Sn�)(`��+�8{��aR&Pz�x%�h:T�ÏO�
�G89�Ao�L�M������j	�G[x=h�V]h|�^��)�h#0��k��˫c��tǍ<p�ϯ��/%��oKt�a��(@g?>]�d�=�y��"����Z�7,���B�^�Z�?w�
�y���j���3�� �^5���%;�����8g�t�F��97kCO�/�GE������V��B|�U�Y�1���Ǐrq���Fi;X��p���x\z����}���#M���O@C���xŝ�����^��Z5X�a�Y{�u� �e��3� ��bH�4n� ��Dv��kj����O��M�p�.LO�[g���)�Ǡ��ː��!ŮYL�X�[Gf�8>7<�V���$ȍ3ð<.P����Adl�c�r��n7Ol?&RI�c(��|t@װfB�X�dl����H� ,���Z#�,��_,�~��]�ҕ�IU=e^�o/n�{^-�Ỗ�a�y��@�L��:uM��ѣu]��h��%�?	���o{.������vX2���I�
��Ձ��<57o1,���b�hz�%����Fu谟)�l�ƻ˪������܈VSȢ�N�i�x*k? 4^���#�G�������H
�z���;��(e�BA�8~�G�6�m�Y�"�{8n�qZQ� 준d��G$)�Y��Hy�}7.9�FQ�����ʻ~1
*���;�My\c��L3P�,����+���9Nv�
f������Q�N�}�,Nps �E\��*�"����c�R�����ɢ��#��8����@��[�:�L�t�ƪ"j
 *���'�A5v�*�`��5T.A�L�9A�����.��~�!8u1(Ʒ��D"�l�?���x�_2�fX�� ���_� �,��:䣜���۹�t#J'��w�m�p���`nET�,.h�˚�����G�)�˥ι�һ�-դ9_�z����)��.K�@!��=7d���XQy�z���:�=NJ��8��o���7޾`u�	)��4�`rn6���?u=����ŌMn��$����/�a�f������j��j�l2��!��>{ٖO����(���Fֆd�	;�����Ȯ���3
�xր�&��1y����		C�Q��V�D1�c1`�}aS�mm6#�e�z�Rm�g&"Sq�14?��k{垷�U��?������<��Z!m�@㼆{�*�Z��@�kV�� S+iz%}q�D���_����
��=C���-��A��o�X�f0v�<x.'�..�\J{�FN)޼Tf�P�z��N������"{���~��3�O|:��R�iU��D�-��T=ݩ�s�R��B���
n���r���6����g@���E�*o��7�@��eI����T���yM�Q(`x�z��L~Αj���7��F�r���7�l��O��u���\�
pc�z�yi�h�&��&t1���'��;3�X�5#6N�Ć�:w��@[���w�-��y��*�����P�N�S���Ԟ�w &O̰n+��=��#I߷mޏ%��}��R׷A�&(}aK��)簘�KHev��H-���X�Mg�~êY��`��Z'�y����yZFhu�p]���rSR�m_2�J�E���Y)�Ħ���XZ'�~h$��<f���cis�N���Qi_��'pM֩b�[�%��4�j@������O�k��$L�J� !�^�RoK��k�%�:
+�i��/Ŧ�c{��6�\�1����A�����5�$���ҷ��rH��Y�#�{��Bg�E%�::���,��~�c^�x6:���h	��0Գž��g�#%��e�#1��_�$�#��m�����t�*�D�B���tO��|ײ�`�'����"�V���1���#�_���q��:h�T��,"��2�oI���e����zSԖ�wm��^�����c��!j�fN���I�ӝ�k�{�U��+��ࠪ�=^�b��8]���Lj���k�+��f`��h�/���_��h2��c���Z�h�t����r��
�-A���ls�ϏL��f�58o��
�Z���LGY���䊮5�!!���e^�ї�w�u+�g6�3���P�O�gYMR@.Bm��1� ��'��wi'/k�&MMeF�q����9�K(��@[p�k�"p�KN_�,��X�<�^���S1�K���s�G��^�FLlu��f����N�3���Z�j��(n*�%�l�~U��#����j�p`@���v7��~`~^��e=*�8yG�i~EbW�j1����=AR�X-(�l]���,�%r

� ~:����hެj�>�h�8�y�B+������лmJ����&lL|(�����^3f�<��TC�|�k"g�A^ȏ�3�#�׾�.?<��Hs>5���9���X`�~�G��r����C2Y��/ޟ���L~���؜���`�:z�<�;oD�mz�vݟ.�l���?�D��ʮ��$��L������ó���M�$�)���|��χ�BF�X��8�Bi����mU��w��2�=V	�"lB�:�H�8�\�*{TJ�z�>p�Z³vW�K����<L�Q�x����(��1��f
�]������5�2dz��@�ȭ�X�0�L%�I�;�/Bm#�ٮ��/|@D��J�Y�"2,4{k�l��~��G���7ɡup"i�Um̀��Y�#m���x�(M�~|j�tX>���K���U��g��x�Uh����M`��4�	�N�1�I�Xi����͔�w�-���������͞Q��g�<5�-�5�*Y���"b��� )���`�[�SQzt)�*)�%ϟ����d�fo����e�ln��*R�ʅ2�c�o.6�X/K���N�ō���q騫�r�u��e/�m/�����fF��[���pH�/�/ʂ�,y��@A����5�����[��'o�ك=����15��?�	�xHݺm�"ߑfeE�i�����i���ݡ�"�c}956�TR���h}`�5k%f1�eG8�s��:U�m�TT�	r�p�o�l����{�Na)��͓RIJ3��S��e6B5�_����J��G8;2M�x��4b��߼�~�\n l;�3e�R�*36��J�2lt�-+�5�U~���E���c��LoP�����|7��&�+�m4��yZ�M
Y�ۿ�u��qꮕ\֮Df"�R-��I2��io+XW��m �;N�L�ԲG�~�3��4�W1oK�~���"N��m����t��M���Ii��&.R-�lO�G\�Y瞥���?�A,a��*�E)A�����"@l��?>Э6 X�\�T�PG �b:*�ZCXh����}V{޼^8N�i�띴p��]���'�&�;�P���O��؀L�	��������ߒ��|0�Q9i�L�����dH'���P^ʤ� ��U�f��hC��cb2��C�[A����;*��ob%p�ϙ�����dX�}_ʾ+�J{�C��jf˨]Ԡ7�TgR�����-n��̧�`F���G!�3c�`�Q�Q�ą�Ҁ"TQl�d�|Ч��z37?~�'`)z�A�DR��6j����ݪ2�ˀ��[���-����KS�
��xS��N��Ww^��T�Z��Su�[|6O��I�p�A�
3#�䔭r�d��P%s����f �(M���Lo�/�:�����K/��k�`IrV��u��a���y�b��r��LX��n�5||���pчz�����Xa��W��wC� �Gu�CH�]�0����3�/�B0��er�'"����H�*��ю��^J�K�Fn��������f<9H���އ�vb$&#@7����o������G��<'��F-�!X���&=�uN��g�q�S(Zc�V�6�C� ��c�*���Ѓ��ĵ-(?MKdR:n[���(wOG�ī�l`$��}]~��cDch�f�r- P��vo���>�[Ȯ�豯8!������+b�!��m.z��Ҝ�R�ר&���j�lw��	S�؅3F��w#�|ak���E8>_�ՂKm(i7�C�� L��\y33g�W����Reɜ����g�������gY"��3�x*�ȥ|����A��>��7�a �4TC|�!:#S1.��"�K2���s�.(r�2n�3?{�u��* B�j��mV��3��N 0P���;7T�Ѧ���p�B��aWe���߼=�ƽ2ƾ��k��OA=���(]��ا�?��6�s_{0IVV"嶇�sr�c����F��>��35$����zJ=P����������Z��XU�}w���K�4;b2}	svR����b�ˎA��wK:�=��4��ǆ<.[j�u<_�� �Q���2�gZv� =���.��j�kRaб�W�X�7"�iX�E.�@�NyM7�W	B�����Q�ϟ���/��1P0�F�V|��3�بE�6�*�a_��.
��71����}!5���̃][���Wa�!�N�k�|����t�Г:#CH��/G��_�3�2V�QjW�&/@��yQ�.&��E�v�����8����H���+�P�殓漂׆�m@�7��}�ҁ�V��$��}%��xc�=���3Y����F譤#�u"Y�����x��`���hBLPi	޳[���7������j>3>���/e�'-� �ב���Dv�H��%c�قY��l$��]��}1��u��J�W�c}��{ p ���t܈���j��5�H��V��>_�'��U�>�����%�M��*�l�χ�m�[/⽑���h���3r�V�Gry��^T�9�	���7E�a�Z��%b�����D	�"+0�ukP�=�Ն��&e
�����33��N�vW�(�5,l���bc����\���8�xa��_Bҽo �P�6$^������o�P�akz���T���1���v�	e�׹�����z�29��q��F�s��Z����}��'fv����qX~�ħ��v���6�ʆO�u�c�7t�� �������#k�f�,����1�{�MG� ��H/�Y��pTWcvl�ߺ��>`��\�l���4OD@m�!��C��t��G����$�crwŧ��u#�>�\���Q�W��6A�юpȕ�W�(2/���k����Ԅ���+��Q�2�`:�4M`���� 6�d�X��O���p\�/�\W5��i����;pJ<��7�y��/����a�R>��4|��DFm����ޜ�.�+G�u��=��]����F_�e�D��?����	V�Ê?qg&�)��=�M(L����S �XPG�I�0�˓e��W^og5Gm�8Of��4>�/�e��1l-7�l��:'���G[��y{���1���xi��Ƭߺ@;�\0��ׯ? �=j�;���B�G�&����㉍VGx$R,�VAk��RҼ��e�ԏ�u���0��"�B>j�A��f�߶.2�c�Pidt���� 8��J�H��c7�sN�Ĩ;�a�\(��߯κ�0v��A�Y��m���t��?�-�AC-u_hLH��K����<6ˬ����RI2�ɼe�!��-:�w
٣�0Xu����pp/8�?_�ay���]���(���C���ݦ�G7��������_$� B��I���d��t����]C~��zY��2W��ux�W�$��.����%uK;�I���0hv���{�;�-����Z�uhI@'ۼ�'���cܛ!�1jd�BV �m{ߨ3�-z���cU{�""�yX�N� x\�U�m+;���S���!�s����$�"����@62K��#��6h�Dh�.��"k0��I�zM1�4B�|0������c��
�c�����C�3G5<����+Wu7�C��e��'�([S�S��JSt4�����>�[�s*�}a�zx����8~�qM��0��!�{��t�9qv�f�q�d�7�t~9Uk�y�RDA�a �����$����'�h�1����I4�jΫ��8�8�qt,19IB��I�؞kHeX}�?��γb�=,w<��&���Q�>0.Yg�6Qø��R�W���IL���E$�~`�r�ɰ�4"���m�C8����*,_Ma���B��*&X��W��Yp��� ����_����Jjy���
��گԍ�l����ҳ�(]�#�(R�e��H���~y�Oٍ0/�o�㏿��>���\}ģ{}�+-��MzȪ��Y��MӔ]������3/5Pf`]��+�ǽBnt0��p�eMl"�b�bW�Pӯn�<ȹ�cKв-j>1��u����k U��1��5������4�	�`*q�Y޾?-$��O,��C��z�z�2?"H��8�[P_�zgӲ�FKGp��SJ(�9}����A6]�-52����9����k��z�������{��t�/#o�=�s�h��t�q�K!|��<��k�eÑ�"�5W9�ڛ����t*��H,�a������	���M"�Nb��lzZ��I��3�s��E��Q��a�8.��F� �
t�0����Ĭ̤+��UB��C�
g�J��\�IU���!��Y[�m��d��5>�
�Z;W��s&�9�t"4ø4I�G"�I|�s�n�f��{J��6�%ܩo��wVg�$w���.��C!0 ��X�pг�q�1�|
��ԁկ��L�g5�*�٭s�L�sud�ܩ
��j��P ��?ϖ���(7��m'�n~56�����X-a�cH��P�,64���d����@�*��vm��W�غ�-�W�Q�i����!������W>��
�&r��ra�i�os�x|�L����2�]"D�����I��գ�$ܲ��ï����6����B����%[���\�)��M��pQ)'����I��4~�'pk��1�*��aK�2�^�2�5N$��=�(Cp��J޽M+&c�d�Զۋmjl�m}Q�T='9}��7�~2R�?)I��(yvw�m{|�ʁ���y�	4��)
����Q(�`���Zkd�c�82�==nSw�Ҫ�Ȥ��tT�t�2*�+��0,Q��(�ss
��A����Scm�R���^����̈́�D��J�-���
������Z�~���IR��Q,η��Dkw><�P�?hT1�}J#p�Sx�����4��}�� G��_���'Q[�E���� 5f^��j�wyڔ���p�|֕�m��6�ԕ�9H�Ȣ�W){�
�5}��?��.��gή�|m)Ku�x��1��M��H	��X�7�K	�=�o����F�0�d�Ѕr�?^�/��.�0T�@3�cn��o:.h�3�1x��6�F�:�ҙY3�=�CQq��޲(�g1Kf�v�b�������Xvᕪ4T4s������]g:#�w6ސۙ�m yT	B~�.���p��D�~��/*��"}��\1D��QAc {��q�-9~�V���%�<� u����ǭ�>��AS������BS���r�	�gh�uSB��Dy|��a�J\�ED.g �g����b��rϾ����^���먻�zp�0���կa��x���x�Ǡ�g�0��F�{��ġcb!*�؊�����;��wQ�;�VLU��Ve�&"f���ԟD����N<�3l��ҩ��?�8A �����t|���-D�M���t�u��pҰHR��Dq��>�(4s$�_�rG�*D�����ds0���N���(�����(�
냟c�������Ҋg�6D:��c�!z�KC��<���\��(��'�dq�U�[fK{�钨yÎ¯���Q�6��H��F�Ep%��b *���n�Kp2o���z�<]Z��0�W!#�]�e0tr���\��#ឫ�vG{z�g���ԣz��z宴�$*�>��������+*+}���4B�P�.���9#���
��4I���K��Z�z�����KK�Hs�b�a� ����{�
�20}:�ϰ����8�ye�x��'��C4&i�č1����-���8��9���(:����m�آ	���)�9K���o��C&ҩmGÇJ��@J���	$]�;2a��a-*l�v'���-}���33�u7�փ���[�<�(U�|sH6�)����c�AN�e
�c��4:�k>GH:D���Ҥ�%88ٿT�����1��+�T�[01��MC�Map������l�������F�Jq�~�U�Ȥ>���;��^MJ_�4M4��T^�+%'<�[�f�)@�d�����M�]x��j����swz2����b�$-���ʉS��K��e�:����@P��U�.GՑ	�RE�AK�Iw����#�����rd����!!��n%7���ٻ�`�=޸�w�o슙e՟��U��%�7D�
!|���v����؛Jz���?kp'�	O�AYx��싹�#���q�6�ۄ�����f�sǘGB��M2}x��as�����=�x��6�J�{���c�~!V�J�;\�\�3���}���c����ʀ�X2�(����9<�~F��vߩ��k&�?2����ᵘ��zL�Ʌ9_�����l�_R�wY�����7NI��4�y!V��!���
D���1D�u
U)}�dr�<{w%��5tUe@�n�2R7��Qw��	N���cҌw[�SR ��9�!1B���Y�
��!ʒVaW��gf5�Q��o+�A�FX^��H����M��XZ���/G�! ,��ax��^��?A���Zve��.�H!:r����5�9��̧�eQ���ϧ�XnЍ����#O�(J�Ql�9l��X^�tf����*9��xwU�|>�1�� ����K��p�7�tz�����
H��~C�/���bV�veBsq��ſ�j$��������ϒT߲`ݻ���׌e,WID�ݾJ��w��GG�/bʮg�P�Na�91��B���a��d3`���}�� 6/ϟ�+�S�Q��ǷPʁ���t��lvF�?����tU��#���)���
�*\;�v�sL7J�	?h���Tn5���Ŵ!���'XZo���sӜ �݌a�)�B�Z~�d���[�´K�M�'��:�Ok��^;�D��f�Q��)��E�E&�Wv�bԺ����E��@^s�z�i}c�сbuF�v�Y�g�_F�8f�, ��Պ�h 6�)_�\�9�#��v��N�"��m�o4�Q2��G�H&_�#�w��H5��o�7!D���;9[̡l0ޠ�1)���ݲ��f����������r�d*k�ƺ �t�m�@L��@=C(��ƵF�������Ô߲�Ls%��M���_��D���`��V��^V!���4��E�/�BtU�%�i5����E]X��k�:�ZAs���5�
!q��	rGJ?�f>_����d��B)�`�9}��<N��u_�PENjN�cz5[yw���!���z�jrV;�4dQ{7���>�
�t�|N���+�1s�V�r��t�C�������`i�J䐉��˸RA�*v��V��u(7���g��Ma�C�-Xł�����ńӱ
���]�y&��M��%��b������Fv�Ω'Sr�=� *hD~� ��a9�e��6�?����>�����
R�T��$&�M���)#�)/];0�(hΨ�{�
ǰn���νۚ8���T���Z�ܨ%`,PT��|��y�R����AJSh>cI[B\^p&��^U4.��%j{��)�������+Lp��
�ؤ�����;Ŏ�7����7���R-���s	�.�`Jyp��':-&-ԯ�I�J ����'f����M������PH4�^\ț�h��ɾ�\QP�h�'[�����0~W`��څ��(�e0u���&���{Së�ze~(� �&�mN�3ϐ� %{Z�I�*L�\V�L	צc�.�tf��-�"պw%4%��	R�} $qN��T��G;���;���Ҡ�T뺏s1J��<�I���G"L��l����KL��:hgb�%E�X��,p-s�QX����]6 	�t���g,��FK{[���ɊHJ������2w���;�<��W$�"B5�{���$� � ���?�^�:X�i��%�&����`� P��6�$J��+j�,5�1������[?wQ�y>��Y6P}�#��-��A�S����+���Fԁn��pcf�������*~�$`Q7��1o01��UU��`m	�@�iO�tZ�)��r�)w��6�1��#	�w&�c��x�b������i7jd�}27±;F�~��]_���٤��4��'DX��H�s�Þ�q5���c�-@�Bկ˓�3�L�M�l��������8�s��uy����/D=aY�{I�9p�Hn]&�?,�W�b�QK.�u�\�HT���%`�-!ӛx�x�>b��X&P�{*��	�����Դ� ���)(��(��s��r.P|�K���;���M�kx)4�w���rڑ�Gr�C,��1����_3&|�����v�ңx��a.T���0� �Ø���s0�=�w:�j�C���2�m�+��S%�z���7� �a�_��M��Շ��;��e���y����6���d���f�.�ߜ�Xx���]	í�����K�HDc"qf�P���28~`�j
Ù�'�|A������b��!�8|Q����;�_PC�`-ϓ/�i�}��3��K����$x��gh*@���uk�Cܠ�1���ogo��W���:ۢP�$��	FvYx�������Y�_����ÚO�F�yt��٫�4J��}�<�̗Bܽ�(�ı<F��=4W�v� �>):�����d&� ��$�z �>Fۧ����D���Ѭ�\q���鉯�N��-��G����&H�#y��x�>f��D�^'�h	˧�q�� �]��٠�N��p��+�-	�G�n��6 ��O��]�����X��W���:���д�h�7I��� �0r0�����iMݽ������f0,#VG$�
k��k�7&MqrIm���n%5e��pe���S&��ݸ��ĝ�@1��X�z<"�b|�Gȶ�0�]$b�-��Ps��MhE�K�Վ{M��ׄ�'�9T�JV�n
�C�B�,���Q�$���r��(�	���X�Ǡ��%��b���9���k*n, k����	���T��m��ûE�Jv��ݍ4hۋ�3�-!8<�\�c�=}&Q6����� ���z��tҊ6�}* \�!"�,(�/�ux)JZ�B2N�<�Y\�e�.`�D��7g
=�s���E	��Ac#[��uK�;�E�\t5�a>��eB]oW�7��{]���C�Kh�P��~
����5�a=jS����5��J��Y&Ÿ=�5������쳪�2�ilF�HNN܄�o��t���?q�1P�x�?�f_=I���Qܓ��#�a��
�h.[��5.{N;���vd���E�C��/Tm���xc��� ���K�4�9�9`_���i�Q�dp�B&!��}�mVv�wV����S��}��}z���W�{3�m���ba���_�c�ة�b�����s��)l�M������^�׸$ͫ�����
���VԪ7�r��8��=�\V�kה�����b��B�/6��2Y�gm	��.A\�̜o��&n�1 �H-lDm�I%DMZ^Q&}�Sý;��=�_k���:�����z�s���bi�#���g�$_ld�_[�T�0P�*���h���`s���i��0c#&PD6�DWXÛ
eK����n���XL�]���0�R���0���w���WZ����?o�1.���0�X�C^�9�x�e憘�U����Ă��)X���x������.ɽG@��y�s_jA�Ш��~\>5���4W.Y!�H�:�u���)��! V��NZ��0`�^ea'N�V�����I�M�
zo���M�#,R���0:����f]��gb�|-��p��J��?�)*m_����($xF�s�() b�)R�~�i�x@�����G�P�����lض���]f���L�,W��B+&^y��L�"����&�B��]{�>dfG>T?��c�����;K+��.�um:6�3�?������b}OC�<!��,�?��.sr�8���{�5q#�
m�ܑ9��;Y�x�K�m�e���v���3{����`2�A�>�4n�=߈Ť�F�8�o���7Am��j���jq�e.7R���[��G�ƿ>�q&��X��@�Q\��z�q���Dk+���^�Lf̰�(3Z�x�s���fVSx�GU�碑���؆Հ�lv�4�_'�I�
R�%T��q��E~,ՠˎd^K�U}��[�0KՋFԓ�G��Z��83���An_��h{�r�k�j�M��P�B\Ez���0T�B��y���~
��j��ϯ���ʚ{Ί^��V�B=zT���|̉�����X��5�'),@Ł*�3@���@�{ޜR��-�St�z��?�R��U:q��ca$
�V�z�3�z%���<��.%����n ta=��3	��U4'��:T�΃4Q���C�PFz(�ؠ8^���+V{�#�V�G�����I���6f�,�'��<+�lqٛ����<�"��[�6���kX��Ru� Y?�|ˇè��5"���Vl��Pf(o �V޼��nOMT#+8iS�	$?�e�G�	ޟ��;�D�=��N�S
�;��W��o�0�s_�K��	K�Ë�l�o�1W�~�����:����ZY��p-�%�1$�ƒ���*.��2�g.��)��	�tׇr\��k1>�P�u�����" {�uϣ�	\�l;����n`s+�Pj�^0O��QPz	:D
�[�1�]d8��9q�[�I�τ�$���I(M̹��C���i�%���_�J��L��G�U*�nX��'�/X��P�������u��Ԙ�W�9���l�I���l�:4<�!��Ƙ�d�t�f�ĸ��	"[w�;�RH��K`�,�s6N�?��*H�_�ΖV���s4�B|g@���j7\Z��(橱Pw]*^n������=�Z�������Lj�~���bx�&�8�����Z{�3���U��珯e�-��x�ⱚ�	�*%6��̷�D�G�q,�ҍ�o�:u��te����(�s�b��S��7��˜W�;�X�9���_�0+˴��t��c��v �*�b��n�Q���O&Є~�>� ���g�Ԭ#�ɺ��e*ʸ�I������rD؛\f�$ԑ]jP q�Xhb �M�0��L���V�2�feF�:����i��y�7f���H�T�!��K��9�=�$�Or�=9�
�����.v4� �W_@_��|=��~q�pGM�o6���q��uΧ9%9!D��P ����j�����+Cr� �ms T϶��yZfVM�rv�F
����5M����1���֫'H��='^B~/N2�>�~��]�lkFg)%a�_ �FLDF���-��cޘ=��6O�׷�B��[d�m�J�6I�~�T-�?���k����J���f��;P���n^�I_��&k��ശ�kz�m���
M�2�,���>���=������E����D"��*A�e�}8�����	1Z��qY�S�V�51zC��Y�'�}'�������F����Nn�ːp�`�RDA�/��]���e|��9şW��5G���D���_�BL��Q4L�╉/��_�_�sT�����|7��cL+�	0��QAE�w�ɾJX oE����*�|�G�$۸i�}=o�Q����8�ޜ�4�~�cU�����k��*�뢪���cfN:�gdRWX�5�zu��nR��X%BV��=-
\���ۓ~�5��K>���{���������z�^���qwV~�'�u��M�8fh+�_M9������l����ɧ=��I���䶑�8.�`Ca�̔W���z�3:IH�����"(�;���XRn�8�z��# ���,6
s3�J%���bxW��?�I�,�j�f�/�wW�,�H�����\��U�|a`�aMa6+�
�{9�����f/�Ÿ��>���P�����b/��;�9��t�ь6�y��E�����縧�x=LT���Y_�I |t�J���BI��l�3�nj4�r=�C�M��<@�(��O��6�ۻ*�,�P��h0@���s��R@&:@OL��y���d�N�q�r��Mo��Ȏ�+�N�"w/q�@Z���*&� ��"c�}S[2��h�
�_��a�ɽA�@�����Cs�_�G�J�ۚ�f���*&	�R�7 ^t������r ms{,���Cۂ�29���Y'�,�i>)T?ӛ|��Z9f�I�W�����jit�A�QKX�"�u�4���#����N�VK)(�x6��t�vr�(+������*�wºJ���䰧:W�A��C(Ͷ0�|��h)A�̴EE��&��p����j�姀�H�O�}[o�1���Z9���ִ}"=[o{��ځ-xP�4	�q�P�~S��<@��[mK��k��=S���؞��%���}��?�L�������DUQSAO�Y.2�ֱ��ǰ�u�0M�V=�� 3�>l�@d��MDkD����K?3�2�
i���agS:$�]v���:����,��z�ܺ���o>�z(W.�bٺ:'���ř)�:fY�7���M=�bP���d�?&"��f�fO������))�;�{�an�,�4b�)4�ǔ_�s{s-�=G��PE ���-V[�+���+�$�����Ab�$_,\Z���m61a0�d����/j#�/���,�L�l�lg�m��ꉪ�ѣp��8����ES���I�8(т*��lV��]p�P�*S+VF�c+�#��$�*�����:H��JlnN�K�;���<��$s��,��λ̲z)wd�q�t��I}dKP�p��	U�U;�+vl�f�j�eŐӎ��]��
2&�|�A�7�9�jy�����g�hE/���eӏ�%Ny�W����Zmz�鯿�5ӫ:]D���D1�����䊛j96�p�"p����$i\'�`�9�`rR��$�?�\�2�����צּ�\�$ua���sV�_�v��Y���
�Zq�UD�����m�nޞ�](U �0�<vt=B����"/���pv��lK&b�od4Ⰹ@ �v�%����/�^%�4Z<D�V/8ƙ�bS̪�'u��Xӛ�\�r�f�y^5G1u��G�Թ0�t��ִ�qg�'�![N����|�=�&�n�:z����Z8[�#��ӻ�s�;�ˎQ0_�uw�_#��q$���|�8�Z���O�4��"A���L�
���(�R��ձ�~k\�:؅����	HiHf1�R]㈋�?_�4��������y��7b���ٵ��l�V��1�&�y�v_s���j;o�.IMB�T�}x�F�̯���7���|տ���/�ۯ���F5�97�~���u��!zѮ�wRu܌��+�_�g[�͘>N/��������^
�R\M�zQ�Xe �M\Qd��h�H
S��K���((c�DKv��6�BF�n�i{���j��A?{����9?]p`[+,s��U���j�c�OA�v���İ˽��5���R�o׻��gV��#�����|�<`��_`��Ϭ�b
8����rA�Ep��bKQP����C졹Q=Dd��#,H�֌��kkg�����	P�@qZ̽�^P3�S����G�~�&!nE��6�s��Eīp���nIe���N�%��Uz��d�#%�TU���l������|dF2�at)�
֭�Y�I_�0鴼5`����Ȉ���Ѣ�x�s1��6U�
U6{Cr���9����׷x��c�~��`�E��3�n�7�M�5����Mmm���p�$	_9�9�"�4�%a.��y������*P�������U -���E��%����b+nB1hH8۾��U��"<>����ƑP�8EMĊ���+��D.�-S���?R�%�����~U������I(	�Mъu�l-%��>¡�G�7�`u������g��,1����A�2��4�U�d�Q벓�� _RJ����3h� ��V�ߊE��d�Y!Аs�)��\��@�*�񝑰Hv<��h$�]W���z�%�H��.% �	�)Jޭ���6��u�F�:@��Ŗ8������w��zJ�Rv��l�;6�����l�`��[�$s��]o7'��'[��q������HBf��A���|e� Î������ٶ{w�#9˙F
G�CU��5!���O摑K��e<��e�[N�5;�a�rj�k܄�1�n�  8�N�6+_	���D)+eܙk�od�@pB��_^%�V��&����K<٘Z[���q���}ܜ��X���Az{}f�>�����A�ج-���I]����Y�i�^W.�����1�h�>�
���#��2���3Lf���X'SV�a�3��/E^�9�O������!`��?C:��]�����[8J2\�
h/c�i9�P��$�`\��\Cm��j}�C��Q�6��hQ�@�{&0)�a��	f����/4���d<M��)�(9}m�s�&�'UvJ�����rD[`���uW������ ��l�3�2iN�>�+��3L�>YS�"-��Oý��$K�g�vF���1gDG�k])��*�&+��$�i	��GT��>�U[��!�Ǒ�����o�ΐЌe��R���H��L��B��vM[yŹ� ǻ@�9��wת֋��DO�IO��4*evr��x<�Z�3Ɖ�r�=��o��(�����>�C�{;�����e�����ʈ��^���;�آN:1W�
�>���q�������+��u�@�DRtבfjzp'�P�t���m���<7Ieߧz��*�/n|�����q�tF^��e�S���W�I��卬��<�r_�2UeWs03|����4�Iv�]>e^�����CN}U��v�L�*m6�eݧB�L�"uHi45Ufm]Y�ZB����a�Q�cd<h����/p.N�v�nVMi,�^��_��.��RN��#�J��T�`�	I���EW/c�+ C
}?V��zS����?,���v��1K��9��UwZ�F;5Q�Y�|�tf��r�P{�jOq��C���s�_2*}g�	?\#o�T5�~�w��H����1��Y���c$�X:�j8�]��m��&Qh%}}�w����`�l�%{Xa%���\VZ��!d��چd�Ï����,������\:/+1���P�1FF ���/��aE�ofl��F����L#���q���K�!�(����z��.�θ\+��;Ag��i���=5���ﯞ��A�N��^'�Zܠ�u|kO��J��Y߽�z��Q�T��C}�����P1W�kG�D��9dձ?/�򡩺&�\l�:�3It������X�����'�(��b�iӥ�{Ds���v$��/��'>�J���LQĿ�9HT��ϔ޶������{nɄ�35L�:�#�$z���S�T�X�y�l�͕�81���*W���(��B����3�5����=�έ�q������g�pɣ��pe��WH���mLAi5�7V�.�
Gi�DM�����t�\2��,�p�T��(=V��s5^BW�T �~���o\���K�L! p��<�����rq@jh3���+GD�V�+
��w1AC�XZ?Dфk[E��������X顈ZA����Z�+t$pG
H����#��S;n�"j]Tl���z� �쥸�Шv���O,�VK����$KA�?ra^�у!p Q���ڤ���wI��0��c;�m]��Tj�;!�6��	���P	<.��C�t��y�h�&OE�ί㊙i�� sn���9 -k�o��mP���<�����������Rfc��CRk�����¯j����SXߚ�>eQL�54-П�Veq�!���*���r�����ӧ6���I������L�멣�y�]���) �h�
����U��z���Uth&��l��9��J�}�9ӣ|M�˺��'t ����\ ���9�Z�b1��U�	�X׮�+)�Bs�@2||�A�:!�|`Ã���I���[�N�p٢��]n^E���{V������,$�g�uFu��qwm�����VR���U�飇m0M��b"�(�.x��nzK���b\�uB�~/�a\��:�$�l��F���
ËK���
SZ���cW�@��lk�)1:p�I0�@Y��re@l��i�2��C/��J������`�����u攮\c�mi �p�S���{�����ZЮ{q	�;P��,7V��4o�%z  m�ߎ����(�CZ���Jv��r�*v4��Iy�2�ׂj;fJ��Y`�EݗO���lD�A�𬌷H��.�Oکk\X���ʌ���Cq�i��@���]�Uv��D��`�*��Z �O�����(	��!�.J5�V���� �v����D�`f2�^䱷0^(|�b�Y�̫����}�5+�m���]8TɌ�~���d�	����UP�>F��]���!�x��w"��)�����Aw��e5 ��~]�i�zi�~��K��E|�R-�រ߭HrGa��[5�lR�$W�1�Gg�������:!ؐ��Z!�S�m�.B8��d-V����*�_�?�*7#��c�B4�]��6�+��"|�w}uK(���6��x �x���3U^]Nq��9w���nQ���&m&J�Q�|�0�Dñ��Ɲ�*����s��u'�N)���Xu=�+a �Jd�7���,gSbń+ĳ���W���>��Wj^|w[��r����m�_��,���b�`.��G�Jp���qA�}U��o6��U�/����'���S�:@�]B�������29��֩m�f/:��W����!ПhB��z��Lg9?�޿�G5p��<]��&�\�|�c����5"�>�K�ax��c���j�N�syu�w���Ӡ�p8n��� �3�������wBŇ�ꌬ��!⤇o_��e�5��y�D��&�����k2�2�3x�}eds�/�gړ}�|e�{�.����I].
F��ڙ�J"x�E/I�?$�{*�|��k,Bb���+�
Ѹ���vF����ol	l+�����ؽd��B����-�"����{� �t��#yT$v�V��]Q%�$�G��*D�x
N	A�O��eM��<���o�!5��)�������b���Y��Kvl���}�jd��>i�qMŐi�qp����� ��ҵÈ�4^�i��L�U�����%���$Ɉ�N��8��"�Ѯ��Bɛ�f�"�V��O*=��}���L���g�G�<��][~�d�׎�G���1��<��!���Z\(7�@�Ncl�on�h�e�C����_�w�;�Q��$R����2�+�P$�;j�5�\�7h�a��q��1K{�e�d��=#�Y�dW&Y�D
���b�u�\�'�j:�%�4��.DrG�A�*�P�BoÜ7f�×���Kj.cr�ߔ�G�I��A����f����_�_"$�p��_��1�b�R
I;��vF��ݸÌt�{V�A����;d'lS�2Dmi�����EOD�1^���l�
�(�ILڹ��SEO/�t\�A��o�4e2�$�`:�;�b����w�CO���&���N���i�g�x�*,�ൺ��� �U���̦��ܻ^���%D��R�3�.T|/���A��%
��	Uݼ+}s�Ӷ��@90���fH�_�p�jh{���ם�p3�wuW�mr��'~ 8��[�v�)�����4:��98���*�D���N��f.�r3���ܡ�t�Z����.D&/Um����.]'�8!$��J�}:u�Ӝx6.+n�z"IUCz������o�C������0�Kߙ@}��"T0�y[�aV)%@���C�� g�����@��B`�s8�~�@����3i'���=֩y�}8�bJ�9_J�I��3�f9�� E��h�M4-��;Ykc�	Hg�um`@-�*�@ D쟉ڗ7�G ]��KԊjC�Sg5`�'!M��Mw$}ڦf�i�h�f-U�tDHM񾓰#��>Qh���r9tg�Y9� Tf�*����"���~L���d���޳��ӯ�玈�yQ�"6� �t�87D�_g�o%vP~߿������F���c���ݞV75I�aڣ1�v���G!+�y�3�ƭ���C�+��Fqzkql�'��cC��*������ep�&_:�c�C�X��<Ž�W��� �cB�&�V^{v�xIG�9������)!���"h� �)�c!�H�!J�u�$� k�y�o5��Y�Ö	��W������X�q�3�J?/[v��R�A�`��#�^c�q���K��A+{wlB�L���'���J'z]?G	��>��8.�(&�U+���S���2�I*өL��ɝ��+�Z��nۧ��!�^��Gh����_!o�z�;�9� P�LJB�4��ws9
%Vׄ�	���F���)��M���Qt��#��.��*��N}ອ4���ʐ�dˑɈ)�
(����t��-EO���4�І��WB���U�¨l��D0r]�����[5��]��Cc"Y�m���d
i$7�@��w��?[��8�R��J�6��2�J���'0^�{u��܅\#������Y�[ ��D�/?8?�[������U[W&�s�J�����R�l���7��ʑp���p)�}��]"LA�ȗK��c0�CD��2`~L�TM�+?M1�<��04��[�-�8ްӹN!L�m]xz�d��܃vk���
��j_�J]���GP�����K�b1�˵W_@�{	q0���oh�=p�TƐ��%vC�WE�@���%�b|ű!�
I6~h�`?� �u��d��/.g�����	�=�u��� j��%o�������5oaBv
�Q�~�r�0j�?D{���T����ԋ]�cl���B�\�1�n$�!u�[�AWl2M�3E�,}Ŏ@[���0�ǿ����%בՕa��j���Ț�2�}l�\��[,t���jCZ�3̈Y��}1�4�1�x�vW�p�1S�C�]��wtG���w¬�L}i����% 	֪ޜPf�r^R���j�hB	1�wW�{���{G��;�2I*�/��,R)�F�ڳ������j��ұ[g�1d���1�z�*�oX/0h{��W]�`\�v��=�f�7
 k�J̓����p1#D	*AV������LU������fW�[�۰RbRZ�<r��"Sl�� ?<VZ�XL�������$Gh�[Mҙal�ȿ$�m<����� \���9�ϕC`�_���:}eܻ?F�{a�I��*��Є��ܨP��Ţ���{�z��>��V|~[%�a���Y�ц
8X=q#��ˉ�RpJ���}��!|5M��_i~c{0��%����n-]���,�D4]+�Ng�S�o	A�x�7���v��nNI�Tdk��+��P +O��o�!֧��E&4�T���O�̷�GCUC��x����n;���p�
4�O8�V袟��� ?�V��gK���%� �D����3>Ǝ؍�P�X�L0��A\��
�&9!����T\��7����[�1�9+2§�X�(�Bx!��^/w?�����  >*D�k-z ��-�,+J�IЗw�#LF�V*��	��z�Y��؝� �+12l
�x�;l�#��{^ߦ$�㨪� YScU�as$�<��9r����t�Y��rghT�L��O�H�X�C���E@�$B:q<���Ɋ?
L��g���{n�����k�v�Q�N�!�l�>E>�fry2��X��Ԯ�L��(� �O�ـx{�	:�JE�䘛�{���gLR�
�c�M��~�S���Eh��%�!��˼ ڨ���E����5v
��6�%�R�̬�bz��t`�I�\���Q����z��aa�����Գ*"&�H���=Q7% B ֕z���a�ދ�`��&��9���C���}RC�x_���j��ׯ�T���h��1(T����'N*�9T�����"	a�X�4�$lL
�其��e��T�	�i�vb
Ԟ�)6)����P��
��k1.���h���v���7i����T�ʯYg������O�S��tݝ�ʭ
���5F���}.|�ViKd��%	��=�bK��)����A�TW��he�1kh|�qiON�{���<������[���i	�¢t�K������ʷ�2t:�80͠I��S��=�T�44��l�h�FZ1I�U��p���^�w�ry��a����H��[��Q�!�)����z��f<�4���H�:;q��ߍG��a��k�k��<�T�s��֖�l&�4��8 ����~�n�~�Dh:}4�M�$�hC%�Ļ,G��u9��.m �5��^T����-񠵽+��A�9h�];;���3=DS�t�*wMZɺS��-Z5�o�@
ʌ������^��=F�T�n�Šo_؇����6�[�����JC8�߽�VQ0��7�P��@�z;(�2�A�Vu�]QM0�?*�`����pI�i؈� ��Oz�`�RU����U>����7Q���)j��lװ�T^�?bj�����Q���+��8�z���]�]dX�����*�G�N�y��J� 53�@z�,��Hz�E§p4<�X0�؏6��:��`�z�<�a����Q��/�	��E @f�:���Op��c�//<L���<C<H�=�|d�ٹ��x����D�i+����Ag�&T���c�����D�38RI%����D��H����B9}8J���XX6N��?	_a&$C���R++���t�9�"���H�����~�{?�~B��YWnPeڻJ4!͗K��} I8GO�X9(���W�����l�������X1���շw"���YN�2���{���H>�w��VlX�n{j���c�6�C����0H���-�jh�&꼥&��V3�պu��\����gQ�d8�&�7_�8����z� 嗀������Q����]@�����hr7���"�͞s,g\�����F~�r��Ֆx9Dh�k4V��)�� �d18���_?�J�5t���%�=�堸�@�\.��j�"�dXEI`�%���Ut�Xf=���0i�As4�t��ei�+}�U��L�(#��7i�a��9�Uo)В
n�CM����p�Sd,��7�vS�f#?�M��%@���l4[���:UZZ�a2�eS�9�c
��a��7x!�[��\~C�����b��3�^sK2L������D)��Y��7�>K� tg���o8��S$�_�q��[:�Jn	��',s��Z����eOn�X���rX�ڧ<�ք��	g!����'����Q��6���r��(�_�I4�D�v��J���B�,v����O{Zw�k����@uX(6��D���/8,��_ǝ��3wNP�[��,P�+�!�TB��W�2�@���AO[��.�ϲm��4��ag�>f�Cwe.�	�Ūs.^~R�8Q{��8�zU�}b/2���	��S�" ��>x&���,	��ُwb�v_�Ɗ����V�U��o��5=�����1�p�a����pAO�l��Jw���蕁N+�LG(�1�ۖ�����b��1��~�ϕ�^������ M��π����}U�T@�S�h�t��U�U!����7bw@����0�=�~i_��������D�� ��/޲��B%*�x���/0`
�o@�8�h� ��8o2ɪF���H�n�t]X`���9i��ik�ӭ��u���k"t�`�d�ˬ�1-��\��B���l��z�TU�yv�旄�zWS�P5fE`��V�k�"�f�60w�\�D�FX�}ݮ=�?)^�=F<��z4/<�s
��.b��p q��L�(d��ƌ}���Pd��ICw��7q�S�^��Zk�%�p!7�{��n�f]�΢~�[����4q��x�h���*h�50BT��tC��VW�ACq��I�Z�9����G/)8?h�%�萸|�"~���IA��dOn��Ȳc��y6���b7��1��j�`tN��{��Z%ޡ
�K�Fs�I�|i��.���mNE����I� ���p�OMD����n?}��ȕ���Ԡ@�fY$��l�,4$b������q�u}�S�ӮlM0W�TW�}��ɝ��h��	x�ϧ�̈с��[�K�C���V�2��ܮ{Ƀ����4~%�26�v��y��{p�6u���=���>9j6xH�0�坟������|[���%�ss���T��ω�'� ��ʏ���9�<���V��o����^0~��s�Q�Y��rķPn�ad2�x��	�O���9\U��y �������Iܰ��_w�jн���!Xy�E�2����҂�ܮG��X���cJ�ص��¶Ǯ���Ǜ}̑�t_^1�[����:)w�j�ۿ5@��~A�?�#w�fp�(���
�G�M$�3����5�P#��h����osX�
�N���	��\ �TA��SF�	N=��$�b��� �r~o�dF�n�Q͵��3��)���<������nz抒�o���!����&�Tr�@��dXڷ00�1�*�,��R<���$��"$^�%;�Nx�������3���xɊ¤�ϼ�yXT��nL�	�,Õ���m$�~�
� XG�-#�9�>͌�����΋Yt[��.j�h�.t�8B#�p*g�����AcJ\�0,u��,�rf�nd��es����T~���"�}/cFO:���L��$ f�W���v�T��<�# ?��ã�T�]4�J��������D���k� mPc,��`-=���a�g.�����O���ծC��Va�qx�V����
~7p'@� yQm��}I�ߥ�g�|U���N�טּ�����qj</�חk�"�~���h`(��`RFT��b&�ձ. �M��]�3�ѓ��s�BK%T��}i�b���pqܟ6�ᾃ ��k�z�aA�����{�7I�64�F���p�2	����(덬�\���R��H�B�OU���C�v������TO���LBY98�pO�f)��,��&�B^&�����{�LF�&_uV��tk96tsD�>�;%P�D6�v��{v��A	��+�����q��{��<�Y�
��r�1�@���4LeWA��e�k��?U*{�� ���D�P�P���Z0K��T0�Ms*��ߥ����;���Kz� �_�YJ/�?����<��Ah�H�&�V]ڝ%�G6��v��]�|���n�oF���q��?��Z8�	n�� nF����򔢏>5-
#I���R��F��E٥R������B���^xeTC��|�v�/%�vt��d;���ԓd�'�JI�r���W��F�]�C����$ڛ���&�+T"M�-�(ޔ� �v���b�geYC��si�����R���l	�Q^�,� �����"�Ѓ����`�\Y�S�ZX���Ɋ�mR�׼Y�#L��v��!0bK��2���pa���3 ��]ǩD;�<{�����K���`o�Zxx�r�����f̨���ʽ!�}��w'��v�2�P�+��T�Bk�&rȌ�m����K�J;)��k���
���f�
*�e��w�kpY�պ['$F]iם˽��Z�|����$0}� �F�V(��S�G�ߠ���)묢����Z�q=�x�	�q+6l�9�Ey���2�D�iq�2�;�%v�
�7Ap2P���-Aut��:�2~����OA��f�R��	)K�w��{y��S{�^`H���ʳ��:!N<��2��㚩D,\iQ�ot��R%����J�EQ�"jl��F�ٻ�]����>��X*�U�Ъ�y��gj 9��R��༃>ͩ}���_����$��6�(|��Ш��y$|�"�j����	w�ʠ�Е��l8�o�`�wc�D���^����~c������_�B�	�9Q��eT�P�.��7���i�6���8"�eD׈����R�v�1T������I����#����o̬VE�g3Q�"N~�zr�d/K�)0zJ�&��ž�� �;!��}H\���9y5#�W=��
|��[�X���e�����׷5Y�؀e���>@E�buTa{)�1����G��?CO59���`�ja��W�5T?�x�a#J������h~UEɅ5����|��z��eu0���-��LnF���|:� �Ꮁ���Mq7�#J gu��@����6JM����/ò��U�&�nfl��@�����>���_��k��K�H$��Lǲdl�j����X��sS�%u��B�Ne����Cx_�T[�e���ꡉ!�����90V�o�(��,��;x��ÿG�܂�O�l��3��-iB$ȷ��'�#70�-E5�B�Z������m��_�H��ۓe':n���2 �>�:j�I1X�~����~$�d ���������F,y$�[�eC�=ƛrY���#%��o��,�-���L�����f~k��d�d����UN|�ӹ&&���zz
� Q��2b���������_r���Cw�BT�J�nǪ��!T
�l�D��|�!��{�u�S�y����*[⳦�jlѥ��Q���U�����tAյ����K�ܠb
��wy�ݣ�&��
R�t��T�Wy� ΢`X�TM����:<p���ecG����]CX�!��Ln-��<S�ƪKC%��2jXإ\8.��F7u�l��E"1�o��0M2F����eP,�%��5)���pH�N�j)T^��Y#��x���H�E8����~�}��K�t���>#z�}[\&)͒lTd`�9B�f���e���R�(�#�ye�%b�|���(�l�\vk#�p�7���!�)���?���k�O	�;���*O "A���6x-�c�Hs4k�_��3��5�	NVV���o��<A*����/[3�Dw:փ���Dl��I�a�q3����}��?�Բ�J�ܴ��*pו���L�v��x\�t�BPAK�(L2��JqJI�NT�#�6��82/2��j��:g�R�3�D�-���R��a$ڲ�"��7�3J4՚e��yZ� �G��@D�;^6Ag�ԧ���$�����1�v�猝O���繫��5��-��P)���
�W؂g� ��'���Zl�I�썷�(�k�/?�>�|��$���z��>�p�G�_
w͔��O�k���$2df\��D�@�$�w[�N�,Fe-��{*9���J�~�u�V������z��.Ke��PKJ�	h;޴�Ӹ)�0���#�(��q��� ���!:zLiK���'k�eTB�m���h	�i�(�'�
�T����4�}��c��y��+�/�X��^���JM�����2A��S/��O��vs�у΢���fKV8L��R΅�t���j'���N���;�����C�ؘ����s|s�U^���k�B���ʜqƮC]b��r�T7�� zr�{@&M�ɤ�u$o�1TӸ. ��|����]8U�[�PVS�m��2�y���p:*�1�Q8��##�����{{�7����ؑ����R�O�t�Ej�=���cZl��Cah���RM���,���cx��[nT��l1��%�hW��E�V �Օ�E��e�[ث�y,�kj�Z
��&���0@ ���#J�%��ս��1>Е�b��ܼZ���0:}s�6�v��f����(�c%�h%��	9�oO�i�� �Q
�?�tSL�F�A�6��0<Z��~���߇n��t��AAz�����d �����Ts���>)�i����s0�N����׷6C;ωl���߻գ�&�,g��om�Di� ��76��������4Zj�zy��/�����Zd��D ��X�,}gȳ�Q;�F�!|���cPei��5u
���~k365k!mBX �7�W�
y#��_����J�� ������������2y׃H�ɐĚ;nqKH�����n��
�Κ�"�5'�9]�kz�Ҭ�`�l���O8��_��5_�K/^oN�銃S�_ZC	�`�F`�Z�xiLQ�7�p���y��-���4=A���o�����6�Jtd��5j�R����Yi�xAsU>�o�/A��#�S����kK78����5�TM��L��!V�_���G����R�$���"����X��l�F؁��zE�Mv�<FB��x��#�����m����N0�&�)QK��r���QN�����E���*|�X1�4�SM���>.�+7� ?�� z���2ʭ!�������M2~55��,?����cO�׻�P�)�Ϟ��[�,n��� �Q������?��;+���k��c��x`Fa&���)��</W��rV�9�% ��B�&��eТk�Kr[�M���E��t5t��3�O���#�3��4Us�
����1_�C���ղd��f+o����e�_�B�)D�����Q̝O�KG�e�x��M���\^͋n!+r��ڹ!�;D�#���!R0��;�>~��*JT��H���d���fI�75�̥�I��a���xF��X ��ї�Q��rN��E���I�*�'>�}T)�%���X��q�Q����~�!�u����ێ�u7��aM�Њ�c>'�fq�L͏�@��-����A���m��"]̗j#f5���g٪P�Q��ؖ�=)�C$�St�0��4�{ߥa�$#�)tV���Q�Q�Z�k��uJ�&YJ��\J������ʃt�?4EG�n�S ��:5`3	_lΌ�J*K��|H��w5ǈ���n'��/��J�o�͇J��K�)UkT�F݇s �3ҷ��,_(�4�� �G�G�A�v�6�|nJ-�����l�(6������T�����b��Ka5��Zԡ8$��!�3ċ�2��ey,Rd��F�h�q��k��)՝��,#!~+���]F4��V��wr�ۢ�]Mt1��:a-KK��^[A�u��X���%�:~�e�q��nM��4�)��F�!�=&�֡�R���J���5�$?��B��C[��:7���(n��B���k[#q����,%^7C϶}onA�����(�!	���-5n��r>X^�"����K�d�R�	����g��R+ޡ$&��0k����jg�>�fQ�TIB��S���3�؆��w����c�f��uɛ9�dG�k9l����7�Z4��"������U�t�NS���"@S@�q&-E�jPnp!1�������TK�/�_�
�z1X�sZ�{���f�ʧ^{��_�㠺WK3�6D~���6����FK�Q�K���H6�45�-���H��2Y�Q48�D�����c[�U�Ԃ��<^��G���fqw�Ǒ��	$�@��k�D$ZqLw��y��VC�"��'�H,e�����H���t���C�|FPQ�$���"*gc4FÀ	�NC|��WU�U� �Vr�fkP9�C�T���r�g���l�э~kȪ�X����؟�q�ygkȓ�gg��&������ ��~�rȇ ��6�bl�o� �Յ��v��[#�3��n@�/.������gޯ-3�ef��CQ�/hh�Qb6�45镴�t�v	��)/��È���|�(��u�s�L�������K��9����W�~��L�3$	��4*����kNҨь�c;!�M�yZ�A�Z�g(D�}1��@^�|�f��J~��v)Hf��ӟtU�xN<�Ѿ��~l}r�_%�`PTR���[Z^��Ż�����%fٓ�D��~��ʧ�W�ֈ�r�K4��'���mφm���g�Y�a�8g.X�l��;�i�>B��SІ���dQ�);���32w-�Jv=�	V���I�'lh8yؼ��8��5$[��[���J�TC���rv�O�����_�6{]��*�!	�ZҎg@���h;�dZ���h0QP�Ո�6^A�Е�y�*!Qp���W&�X�����[g���׹L�*�l&ox�����bV��!�U�8R<vq��=�.�LI�Ӷ��u���J�ն���Z�*sx��n��?np�{��˄�M��¹S���`^!A�m�{r�~�G	�N(˶z�ȉkm>��]S�M���ä�O5 �|�L���\KQC����0���W�4�����Ӛ~�&KXX9�����!%K݂��4��
=� ��"����~����z��J����X@�U����	���ҁ�L>�E��e�_�K�=����0Ω�IG����Z��Ľ����@���U�v���^�p|^J�����]n�����@�����*$�S�*�ֳz8��n�>�t�GPu�քFBCa��a�'z����ۻ�$;���o�)�6���!i�&��*��PpwhToJ��#� ɂ̭�9q���$LL���#.��]<�'��/|_;-��A�V��Y<���Y��2h�[A��1��^Uxz�ӡ �*�X����<cӆ6��fI!ui����ߑYE�m\�Y	�/�ɗ���X��;b�l��SP[EK�/��5�9c6AZ�%/V�)��~��M?��W|C�g����g��@�u_HD[�]x��41[ះoN6/v޹��|+��N��v^S�Q�RyXu�z���Gy�@���\�Y=��Q�9Cq�N�����v�UL�-,�^r�z�G^�{�Vp��n�ح�����"����!�c��
�m���o���9�E���?���W�4�P�?��`�!��'��$zk6���!�������}I�ݳq�71�۶/����6A�_���O��w� ٺ�d����×��c �wǍ�đ$(�s{�9S��@!C�ʥ�w��)�����_r����Vt�F�P�||�24�Ҫ�R�"��p|B��(�J.�O"����+B�ŷ��R��;m������.t�t��9�R��R�;m�*BO0�T�@b���a�M*�]=�(�@Ұ�}L��]@��ʄ��kRٍ�ò����Q����bV&	A �f��9��Ҵ6�+���x������5E�#�D����" ���0e΄�8�oױ�� �hz�C�^�L�sA'���|�U��hZ�WK
�<m/�{�DK�'p�*��T�[�Լ}윭��X�i�I���s)�;��"��Xl���Ch\�q��6�r�Q��JT\R����^�ޛ�X��U�e`ʽDҌ�"z�a��0�>m��Rl�w�"�Z��/��ڇb��cG^���.qRn����-��"t�EIj�m�
#3IT�M�w{$�PL����UPj'�2�����7Kw��.���W���Do�/n`x���f�S&}�+�U<�x�z`�1fm��L�����ׄ��� �e��^rc,�zh8�N2M��WI>2���[¥㾢Q�:Z#���bs%`���`zaL�=��r�D��4�mGI��\�2����9'��Vr%Ԉ%s���h���K��)�DGŻ��������d���f?��R��N�æ���h �ˉ��|8��e�Y
��n �����Uo�ߧĪN��}�n�=�6 a-QC1���R3�E��3��nN/WuӏF����-�?r��#��A�o�l �{�	�>W�$��ګ�vv-������/obd:
E��*^����,>�Fr|�cO I1&@f��x����
)ݡ_����@���(��~�ꋱU����;�cLkuD����:�,5�r�H�X�A�%Y��%lM����
J0[��
���V����B#�j��S�x0�����v
򄣪2��<pp�@w��[BT���6
t6O�;�A�1�j��$�n��C�hz��V$W����p�6g��+�^{�E���4���{8		I�)(�Zny�ͺ�%M8�������6���ךp$wW-�q!a�-����tdi�� KE�+�&��d/�t��`q���?�B���S��H��C���B��/;K�A���- I�;��7+����OB���!,E�9y���nk�׹]g�����9�ʸ���+�	O�+��{���Y�s�&�ڷ[B�gwu�U��,�� k��9���h0F��С�-���d�@�J�����I ~�Ƹa+�����bH����͆�W#��tJ.�E�.=b,�h��{&�X ���F��]F��p�����!!.b�ʶ7︔M]U,?\E`�fk����>#}2��=e�2>�P���W����gҙ�ی
o]��T�-��A<4Tq�A���TG�C?е����q�J"q�i��n��D���<ý���[ ��;S�;��k��H�7����tr���N<!ε���a�zDcČ7}���:��B�)���]�����e�NN���gm��m��"I��W�֧ ��w4El<ĝ�5i���X˽�����3/����Z�sL}�YX�
L0�U�N�F^�5�E�!zg�����ݥ�M_}~b"���/,!"�S�Q��E�^q�-����(ǂ}ei�X�c7�\�h�+�k��3��M�<��0
�;�v�|ݧa��m�;{\�;)~��^%r�i��)�I���/��x$|���{�>{��ќ��͘�E+N������~(���ES"/- ��!J��>���nֶV.Nx��*R�_֥��a���<��=Q��Z�I�˧A�+��h�{r�S��m�nևڊ\�Co�Dyҫ�'���l=�ƺdwd���xI�m��6�K;�#E?���1~�<Yc>��V8�pCS�o�?���.3Ru�A�qN�=��O%>�HM�-qb�!C?��L�]���;�,�������2C�C�Lw4p{h'rs�{P��:ٙ���a	����T�z�,{oS�b���x����}x�F�I�ܐ�T]5�8�%�z[58#��%8R��j� a�^���݈^qK�w����U��՘�DZ+����6�t/������.��	#�8 <�;#�f����4%g5�q0Md?�H�YU�$L*��OI�3`;���Zj;nDV� 1kF�@��j��3�%���_٦��o�� |o�qD�q��oX������H���i���$,K���^
c�+��F��1�M���L�����X��p-�K����?�X �����Jy?	�����m=a��m ��"1�i�(7�b�<�B.�6�����X�C�Q|�b�ά���F�L؟Ο2����\q9D�dZ��w	^�/�[�'\Q:�c}�9]��m�$.D��GV�l^�Pd,�_�������F������;H��>���JH�+�`���I�
�rRʁ%�^˧T �QdR�]4�)�8�CΜ���(�U�pژ�ͼ�@���_1�jZK�7����C3��pɚ�{y��U�z�Z���D���ܝEJ������Nɶ�a�>�n)��>ig�[ybR�� �E5��W��l���Dt3r���;Ird{�j��m�$��)�� e!}��\��w�U�f�� ����Q�ǿ�(�d�/�l�BE�>r��F�]m�|H�F3�@L˶�dgi2��;��m�R����`��W��o;���3�LV�F�:��}����p2�#I3Cϖ���_��>P�����I����ֱ��t�H=q�:���Շ#�Q0yH��I�y%�ȑ�@m�s!��¶D���'������#6B�FW��\�.FM�9;�C~?%��)�ŷ�G�GZ�����nQϨJY�d�@f�sR!���`�e@�o�A;�(����'M��y�# 詍5E��X���-���#��%�d�f��,DgG�&+�a���J۷7e��t;{�W�#_g3O�a�B'��XR��'���hy��8`���E��9W��n�p�K"�L���^#V�NG��(�y��ro��4Hkb�����_�o�'�f2�֡AFa�|i��i�ͩj�1!φ��)p�U�����u��ؾ���$M�N����9����ע�>��It"���`K���-3�Zl�S����sԶa�-��_���g���Pܪ��5o��G�/�PˢP�S��4�^E��a��?L;�u훒������&[�t[�s�_?F�瞍��Q*3��K�g3�t��է�z�(F*|��?�c/�G�t��Y�&����#����X2�uc|}c[h�\ b���'�%5���F���鹳D���ǩC�TS�!=m���V{Z���,��-I�zr*�=�mB��ҫ��U��Q�*�\}�8�Y+J���,�]�	�)��#�0v)�l� ێ��Rd��CS�b�����q����`��z'rJyU+1�	J
�Uw��z�f:�����D�?����7����voi�M/���һ;�Qj�.Ey�� w�]��|}8�^�ņػ#�0Y4? ��8 `��tL�ƺ�OB=���+�ļ�<�=�P��媥UÏ���dE!/8��RE$q��:�z۞��ێ��#ٶ2T���2��>
#�o�M�\�Ȕ�^[�X)�s���N�P[��<���9��=��Ґ��a�y���њ>�p�������I���lߟp�Y��ZZ�B�A��"W���P@q��p=|klH��!��ڻ.|L�W��P�3e7�;y,��r��C�C
se��L���W;6SB�=κ���ɨ����D�?vT�M\iOH���?���I_ ��F�a�}E?��A߃j���\GZ��u�P[�Ov�mD��lTSI\���O����X�64��}�j$?A�#�>�}[W׽ڥ��Eb�l�7&CИbj~2Z���ՙK#�z�(,%�:�gq]�p�>������7k�顇s�޳��w��4��L��@e�Щ��`�{GHD�3���F���! [jKu�أY��g��B1��h�h���E�̲^eV��WHu�{XI7��$w����Wu�zL��� X+Ʋ�`E�K;�J#�`�_ej�v]���{����Ch��d�Շ4��y
�H���)f����0��J�Fx�7%����n>[C��h\���Gƀ!�+���a'&��kn���k4-�ʎ�j{�������GV�=�\��{�B�t��nf$�ƹ�Mu@��Pz%*�33�_�2���-<ҳ� �Y���#�j��%8\�U�A�'`ϵWt�`p��Г�x�vߓ����'����o1+��'�_�/�*0%���QD�*��l�7����VJ�D�o���Ppmo%�Iy-��Г,���	���	�zP��N��p���-�k7����*0-9��{�c4`��K��C���,�`Ǘ�H��q��S�(P��XRbW��|�H�M���b.6���� �jup&_m�D��`ho2E�Kk2�W�o i�p1]4�Dh@�C�k/	�>gF�8����p���<�ATՑ��t�#v(�!�$����e�� ˴#�����@�/�/*q�"UBs�F��o���/��q�S�4|���F0�V^ҍ�"��u!|7R� jVO0j�yOU��������q��UX�C\G�4��t"6�ܬ$�������8y&@u�r$�0�68���B���^�Ϗj����$���w8���J�Z��K-��(�Vl�O�Ԋ�1ǔk|�� ,�F�sΫ��9�1�lԞ��\������Ogûbl-?���F�C2���E����m�V����
��Cp�����\���U�C1���PG�}��_��c_��f3��n����|ke���kA�;����E@�`��O�7Ws���a/wy?.x"�L�}/g��y9f����݂e�Uov��¼&+��WV�F6���7A��I?E�M��6e��%l�Z��*��7NEi��`Lh��p��[X�J\U�*?ǹB���b�F(u0��� �= r��#b�Ж���b���k��7�m:���P�s�~e�eg��Դ�O��L_�	���1�R�'��_@)I|n'}+��`����~�+�~ġ_-����:$1�A�����!�W�T����Y$�䶊a,�Z�Yy�CF �)љ�\F�r?�r�=`�U�q���-]G2�S�5��t#���&[�z7s��z�{Ağ�[FT4Ff������u��0�s�;�N�C��j�#���	��^Oѱ�EN�Zq�6� ��|	�K@ ����# W�d[�o_�z�S�̈́Ia�����'jwլ�LE2��\���1�jn�Z\��̱F��u����"7oOI���}��U6�6͆h�|<��2�`�l�U7	ٌ����&g�e���"�.�����߉Ä�T��T�}�Ԥ`끂z8{Sf"=;��3w �ƌ�9��pM�Kxe����XC��U���*�`#��I����8/c߸L�
�Cv��:r �o���#�ɘg��ʯ\ 7_��І��-0�l��k�-dA�	�T�Fm�K�]���Ty���}qY�@㿠G��AR�)a�l�^��ҙS7��HYIƀS�6d���j�=��a;MOT��)hȆ�ؚ�㽚�YS�.���!y��7މ&��CxA����,O6�. 4���#���`���,gd���\v��n���s�"��l�?"=�FB����'&�����l���tn���T�v�a�+����(� �6�v� ��w��CD�Z��'L���7N��8#I*�����
�2��\�Lb�.�kHp�m���G�A\�ﶁ��WU���!��Ͳ�M���6R��e�-�A�\�W}u;�~��]���ۊ�] ���*N
xd�1��<�����t�*�� �� %��AF�0���lMF<8�����UMӮh3D{%�	r�C,�&ԴL�'��\W��O��ݕ��h��IM�QP�,�L���	��K� �a����y�Π%�<�iU�A@�ÁZ�U��48���i�J��v����t������QDG<!�bP�>�NҖMW��g�D�q~�3P@c��ƶ0�)���e|5���T�jp�Q�B��,�V?J|��������@�qp�����>i��*������$����LH��WEt�r�|���(�|��;��vF��P(�w�p��6-yt�k0��u~(b- ��q8z���y��*qi�DQlS6`L�	L���nf�h����29Ip�a�[�Na�ݳ�w�e�-���f-\��G9�#MC¡�9oTZةP<,��h�/gb�M� 
�+T��j�������=�z��dTN`m0�����L���e����|\b�x���']Z���~�g������e�`�EH��bп�"�V��e1|���bo��	���Q�)y��-���tN	Zk:zq<�m�bm@��!^��EL<�t�M�����-���%A��b�as��B�ﰭ�
�lb]��^���z�֕2p��R����A1v��^4pX4��J�<�*w�P߬(ty��!����
 _�0n�t,�/`a5��_���f� `҂�)3�&|vH�>w?!��3\eFh����F�)��%��x�si7	�w,8����U.�%P*ߚ�4�F�.D�$F��)�]�U�`c��Ⱥv�����c�:���|{V�StA�8~�b���2������s�
/y�Nr]��yrr�RI}��t��a�ޮ0�#���֖�c�2M���d�X���K����	�6v+�-'@8����"2����/�� j�(Q�4�TY7�^��^���ݿs�~�B��D�(�{������K� �SVy�8�J`w����ښQN���"���M�ϙ$)�c��YU��U�|>�W�����P�R��������ժ_�9$�f�-<`�Rdu��#ï��X��s��BQ�d�<��`��tfk��낆H�s��a�Ao����o'/��z�*t���#
�2�*Sq ��Ȇ{�8�����j���֧�"�T@�rI�HI���b��+��l�ޯI�����4����#�����!�����ؗ	c�R��P�i�L�˦W�ȏ ��6��6S�$b<[X��p�l�B��YNX��Q!O����j� =�����P-�]�^�o
N5�M��33Y��Cf�ߧvR��<�����+^i/�����jM�:�9���s�M���֭tU�@1����/X����	��4�c�;	a\wˆ�|ɷ�}6����k�)�3�Ø��~>�Y����阯T���<W[~��@������jN�k�'���jnJ�[�L��{�Y��\��z������jOk'�S��Z⾛>6��Xl"��Su�t��i�pl-�goQ᥂��U�3��P:�r!�s\�;7��;`~�9Zzb[���9�`��(�:QA<3`.�숁�i�M�>������q��=�p���Ps�ޕ�s���j�$?�`�반3�h�3ղ��2�~��'[Y�T����M���-�g�n��+M7�𰾽%p�yE�OD�HdT�t�髮r�a���h���`�9�}q͗t�(��ҽ藊z���ι3��@du--�	M�V�.�US���ޭ%���V�L8b5( Y��Oy�J���+O_E��$7Y������L�UWut5*-�}���]r����k˪g#���U��+�mN�s�V.R}�)ș�}
e�Oy�wq�����ʳ�~[<��ZO]�����fn�.)��a�×�G��������C�*6�3��O6�+�A���Lb_�}�ިE�rM�����iYm�=DD���Ǳ�*���˓����h���Kŗ�%�N~�I#� A�v���M=��w)r��Uv�!m��9�;��R�r6d=���yt2�}х�<3��[.�=g]������`%��,�[�M�C���Z6qO�SHErK�]~�F�����>�3!�7X]z�r�Q7��Y��+�Uw�@4��zYҲ��a�(חz�iT�����t����񛢔	8`X�|�OFo�b; �D�v�m�\�*e�o��OU���B�7�M=��7!Ө�RJO�%���+����j��[�`6'���כȡ�5��P�q-s��tY�v.:�9��T�؊�-H|�A����n��5xH�I��k���F���^Y<�{옙�����$L�~<no��
��͒+���}Y��w���v��	�K6�VQ~׌���٫����|�X1'�p� =aV�,���*5�{��Yˮ��UDp\*�<<�<$e�a6p���n�"M���y�g���k�'�������~(b���fj���C�).8�m�9}�)aS )�a� S�j�ˢ�{�źFAŰ�Ɩ�#˪��M�t$����x5�E�G�`�ئU��^��(]t��=��з�KLYkќ*Շ�����/D�i��ש�F�l�B:�b3�=# �_:��1��x���G�R�˱0�O2x�c�Y."XS�L{fd|���w�W!�-�%��c)�"%2zZt��~���W���SPB4����Bd*ց�]9b��V7_�k	
�E�����on5b\��ʋǜ����L����z��?a�*.f����8 q�MDf��>�nӭ�2}ov�Bn;��b�1듅���ܓ�t�+���R9mVN5Ќ��h�*�	-ѳ�����R�У� ��a,�CJ�@R��O�أ�$�+_3eK�&��������1Gq�$P��S�a5����8���w�n�-��KnZ��][��e0�XT����[�h��p:�73V���`�*���
����j�!��	�{?G���)�������K�=ŵ��܋�
�����	�A�)K�����x�߳ߧ��B�؀�&�*�`<��~����1 ��A�h	�KZI z}2p�x-�}z��>UK��Lf�f��wb�]�z7R�Qz!8e\�{�:�?8�" Q�
p'�ߴhri�:��VxBBH� �;�߰K�C�wE����EOi�9N��De��횸�4�>EJ��K�&���9�s;��!��	Dޥ�B�!��e��l�_�h����72AR�Dش�lV�(2�Kӟ6����d�Q����m��f�/.�۫��+,IVrj���ɗ�62�F�[�N9�͌{���5I�Íz�N���כ�����ַ�d����q�P�?}tb��̌�10�B����T��~޾q��O����i�K��N����J�Y���uX6�<�ͯ�my�)ָg�
�ot�-�(k�K�0GJ�tʷ�ы�Jw�p��3��P�t킷�ڋ�]n/e�����V�ye�M���;8�2�NX�������ӗhZ��w�µ#>�o'^�΀>��{�%IS�5�/9��&A,��Y<���^i���Ǩ�y.53<�Tx�W�	>Le��Ч��r~�n�xă�%Yi�2��
�/����U��SB���=<4#��l9)�"����̱��ы��Gz�xc��n4�Q��9�U"͙�p�aN?%	��b|�+YWUk Ӡ�-5˖�u���T�eMr��*�
�! x�+.�\4A��Q|9�A�X���Y��|���n���܀5�;iW�����*b �Njh]�� �e���ûؔ8Z���9h0�4���#��bMl��ɬF)��I�h;��K!��T��΄χ���tS]8�6��M+c�~M>˻&E$~FX��_s��Vfc2|�(����.ZI�U�ʦ��apH�6�%ʓ�Y�����/�A����k�䕳��= ���Q�g��c��0w&�S)QA��_�$�G��,�̰ �UbV�漜��}לvJG\��6��I�"j��;$(.-�"�t����0����=4���*���T��2�O���0�J��&H�Iꋪ��t�.���OY
�GJ�Wn�ح �������J%M��L�����}k�BZ�ܮ��o�n���Z�,V�n���c��a�Fڹ��&�w�ٻ負�c���-Q]Q�Lky�������ew��훕/�+z*p�)��F�g�P�M��Gl����9>�c���H��5t���4�>5"�J��`�7 oo6@�[4���&���+/A�#p�FA8��^N�oG�1�T2D�������#�2nS�F�ϯ�^�A�'������pTD�?G�Y��� �r��i���N��h�=�����e#65��0g�/?���P��p�#�ǁg�|δ욄�d�钭�y��D-Xb�@w���x4D�������L�n-5�~N�;?]�
y�.W^�MxP6�1���|V��DF��E��G�@��쫘5�F[.�r~��)A~_�Ċ p��P�󬎹��>�'2�%W"�/�N���A�~-Q����V)�k���S�����,�'����(>�'/��NA|6��L�R���t&�T�-�E��P�3�<������#<j��q����W�%9�9�K�nDQ�p�Ke�[R���0��#a�ߍ���9�չ�����S�������*���Ğ�F��� `��:��JX�hD��-�8�! m�.�U��Շ����E��%�}׬��-�m�[����8U#�F�uxc<����;��ߐf�&�s��h��A���g�:I�?B�$�y�{�5��wIȽ.�d�9r��z�����zY�[P��bĚ�92�t�&���RN�ye~���~�ǳ1�q�QQ%+��0��~�姵�L�(L�L帩>���/0`��en��w�a��6�w;p�WoV���;�D�D�T�iH�'���%�r�A��
���,�먐+���cw�W�y�x��VZT�s<\G�՝@A�.uy��w�V��K|�� �y������<��g��Z]�_����*��c������bV��X�MƘ���ݡ�foe�u�P�!�J0!�!���Z\:N#�C��\1Ls��xf�����`����w47�2�O��X�������}�PEO�筵^�>~~�C��_���o�B)�������(��i�EK�TԔ��ʴTYw�貾��u2ɉ���������Ü�H3@`�p5�T͘�x��e�B�����"yژ<��1VߐB�s��L/�6�{>'=�mZ�L�[�����	��(Vº�ӓ(�ص�5�Fȷ��eo�_ќ-����u��c���C�!�H�Pߴ1Ђ��{_�C��p��h�j()�8?[�<�Nu�&� '#߻g@��d������DVv��Lg�"&%&�Pz�a=*�l��ޠwz	�3�Pf�[h"y�����^��J�VR N�Vjn�����V�G�͐��Ľ$ �0��K�b3m�*؎�M�G�0��,C��)��WIع	�������j0R~��A\ ��z��~���QGW�e��'�8��$���є����.}_U2�`�9  qu7�T�e�����+�˾�ٚ�"���0�ZZ�Fr5�H9���xs�#>������`{��WĒʼo���WM��;E���493��*{��u_S�Ap������u�J�����+�/F3[�,H�̑/a	ƺ�^C�n<`�L�����J�L�/
^+�@%��Ўm�d[PK������Ssy��,>�}�15�:��c%����d?q��]�EH��e��ڄ<�8{����$<�z&Q�S�+y�F^�2��vE�:�ͣ��-�3�i�B�B���޵�}�;��ȰnE�ex�������	G^�j��� �;���X�|�۔�z��'�9��
��k�p�E��p&Ȁ��IP�z��0�e(!�U���)b}NYfNl�����n7�h�t�e���`��ېs� |����bӒI(Yi�3pߵ;�y�܎�}#�˔��)�J�y�����ou��$�^D,K��O�i���k�][�j��|ݸ�K?h�	��(�P���2T]�p�}��E���� �sЎ�?b�C�{i~��I����S��NV۷�dI�F�������0C����a�X}LU.v�!DUc�d��pazm�-iC�l�ћ\��z����7i�(��NI�6�kկ{�'���=h����X�$�#7�.�P�RlD��,�a�#P��ӆ/_J|'Sq	�b���gw;]���t7���"���'1b�d���h�3H�6w�5^G����j���o8F����g����>T�xZ�Ʉb2�>]�sX��C�~k��\�Lg-e��w[`�n#����ጸH[_����k4�!��ఛ���J���1+�0?j|1�L��k����G5�B����Ǘ;>��.����p�;��ò�[7�`
�F�Aж0���%����`�Q��?,
Cv�u7�r�)/�d�#�f� q�=�!��k����S4@RFuw!��T�޸z3x�ѕJ���"�-
��s�vȶq���.�RS��U!a`T�.PY��Ec;���{�yFK�Eo^���^s�l�:m��(O����R�jjz�Ŀߨ߬p��b�2(Ecv{�N5|fd&�x�DQ��M͖��[��"ʎ����|����!���b�޹��wJ��;���!t�����7&3����2j�Աt��]�/r7�'�-�P*��w̛��^��-�)N��4,���͍���fQ+ͳ)m��n{c�-�j�!�:�l��r���H"��M�2� �8y�˧L��{� �M�j9c�3����)���)B���N��Q2SNG��Ӳn����mr��u#
��!H>�/eCv/.��t�����WXPYn�^�Nr���-�ڱ���p�:3E����+�pS�9H��b�Y�Ό�x��*<��5�7m�c���S�� u|ndiRݝ�ޠ�!^�K7�F"�oe���������U����j�k��+��/i4��*�G��w���a�~ub���\@��c,qQ�'kTT�l�,�����p8�^��^�@�8�����i�V��2f���ڽ�vSy<ef���h�i�=�VT����vmܧ2q�+z�HX�Q�y P㲽�� �T���u�X�h=,2C��S.]^t�f嶣~���|��λ�� 2N$�����(NkHG����p�W>^;��D��#�ۀ~�f�Et�{�d��z��z5G޼6���E�1��\��
��p�C
� �H��h��B�L����f���h4,ǽ@�-x��y�\��ܲ�U���$�K可���~�F
�⭿3�Q_�¾ ��:��Ğ:�iL�'��X"�%B��:�Y�G�}Xd�m+�L�^���Y�BGS7��Y��p*t���Ay�e�Ȼ�A�h�F�o5���0���	�)�O�;�fX?���g����?9K��^��_���C~�S&Ln�S�
� ���kgn�
I�ͯ�R���K��\X9�'k�^��(��1��I��KD��b}�j�Di>X�WZ�5*I�J
�������	 �>?ݨ�&�[�6�M�Ԅ�?�}l�?_6Ȱ2-�a��Vy�'�W�
%AMe��a�δ���Ue#�.# ��x��v7V�5�F��$��ܘ��D�x��z��e�,�U��u�@^b��8�v��������Q���6�'`~`|,��U�����l��^-��K�iV���w�&�e��'�u�˼�hrPV�� �����Q{��%DV2�e ���ڟ&�)
���c�Y/�Ck��+<���RF�a�E��H�������'z)ۼ�����n�j^ˍ�����4���>�&q�g�*��g��4Z��,��s���"=P�(2�v:�ujx
`��.ā�'�/��^�ts�|!(�_S��UI�u����n��u�,J�aMyh�,���\�1��<�5����L���C<�7��W�LX)��T�;���8��fN[^_�ևs�
j��y������Cx o�_���Z ��g%H�SO0�{_�(�����$�8�H����-m�>�Y~�)�g����q�Y�7����J\#��C��Sp�w�i�f)���_��Y�J~�G�4B����-����B%��<�T i���`%��'�q/��w`��*������gZ� �a�ϔ8(��?�xC^�� ��_��h�'dӋ��� ��c0��|Y�2�N*�Д`k1��<`$�P\�v� J�R�i�! O/��H��B�c�d1���l�ɆT�D�",/y����.b*�/�D���{v��$�[�!� �ʢ�W�&��Sp�"Td�e����&We���9RsI%.m�K��h[g��ϒ����򈬅���ö*<%�9��8�I���7�I��z�kd��=�]#C5�9V���eD�%\'���Pcl�-}�9iY�lY�=1����-�a	�w��TǏJ�Pƺ���������@�R^��?�*��7]�GXC��w��7t�o��'L,fG����$,Z'�h%c������r	*��{�F��I��R�g��iJ4����tR�Ƃ�͍�����÷�4�� (�4Q��;�<	�Q(�p�[�qZ�Z���7O���F�����<m�#N*��j<=�@IF�$ �iݢ�A���!5_��^�e$�Ej�Pm��>�����'y�=6��~�{�tVUe�<��O�g��+mv�/E=��Ҝ<�V�Q?��Siz�2.~^�����&"�{���j�pa�~ @�2�2��8�_�����a�=X���4���{'�&3�>a��6�c�W�j:+q�����B���Y�6�<FM��*@��k^	A�]�4Xr��L`Y Da!X
'X[����N�G+ 0Vޕ�29S�����S8���ƫ-<�K粱,��x����l	Iݿlq�@%H�f���=�zW������L[�!�C����XƎq�L	�k���~;7�C���%ECc�%��C��4�d��Q����������Խ�J��P�����P��ef6Xg4��� �ehl
,�N�� ��-���6�W`�a�ۖ�c��-^��d�F~�3��肠?%���V�;��B�r�]����9�'DR�V3WP�U|#qܚ�ۣ���/.�߈?,96�v-au�푟�U&�h�?f���ط��O�vl���3�{B bKd����������s�ʐ`�7腮`�=�}B ������0c
c	�%^nH�I˗
g��$��M�Ts���ۣ��%�VB�I�i�g�י͘��ʕ� �$xҒ�[��#��ۛ�	��WMy����-��b"�n�N����͙�>Uk��k`6d�^���K�sx[s�C��r[�Ja���H�	���j달��-�:�ϑ���=b|r�K�ԃd�=p�V���
�aA!I芑L���7�{[V8���{ʽ�A�G��A��T���0(�h���5�.=��W�(^d@I.۞ރD��V�%���-��t^Ø��/)��^���IH0�z�M8ԞL0��+�������FG��i��	b��T<b(����bg�����n/p]�������{"��r�Qh�d�W��j��)�)�ˬ�����C����}�%��ӅQr�|�5 ���L��}�N�f�P�z�ŝ��]�Ǿ��L8! 4F��u&S�I�	�������ѱ�܊�i&�����[S�<�f�	�;���d�V��]�n�R���'����U��iQk�����	k��G��).?sΈ�{@ր�.� �&�vx���~��R �giJv�����g{�Ufp;B��,�X����I�v�G�}zP	=�׸��F�E�Ru�=����`��c��6����f~�Չ,�y�叽8J�@�\��D��0�ٕ�NS��A7����h��pd���M�C-sY/�`i0�=T�Zǲ��,�5�Tt��z����BURJ��/	3���)wd�e�7�W��	c$R�����/�Z [\\��6 @�ZRC��T�0azq�<�	�E���l��뤿`)[��E�~i\�P;=�űC�F�ߕ��|U���hM���]�~�/ՙO�Tg���w�ԊY�*����z���T�H�J'�Ē�P�
;��=kH�T�861�4a;p���ջ1�B�g�y��u�ݘ�WĒ��\,j5K��?�VX�4�?�r�TB���3ϺN�efl<�;��Pa��2W���F�iC����1�c#9�X����F��P/�)�5�=�g\<�Rs���J�n%ȴ����˰3ʌ�쌿���y����_b��+Q��Y�@R�Y�M��^O�T{j(˹�����c�u���8h�xFߝJ��@ �a��P-2#�_L�wim����4'����8N͝Y�5��X�UKx�A?_�p�urʪ'�T��ns�`7��:��jS8d�������iV[�v��<�<���rk�b�N���a18Z��ׁ��o5J�^���D�{s�I�焏��'�&���i�D1�fO�p�ݏ�z�ߜͺ6X�p �ݖ���C�@�s��-n�+dH�İ�G@�z�b��%��qQqRtS��[���xo>��bŹ:�
A�Z*���8�}��8�)fVħq��0Gŷ�%����|fx/�F�/�v	VK ��-����Z�ju��	#�P]Y��[��3��F5�$���/��_���[#�\�םϵP_��%��!�I2��O���	E'`/�/�4"ٖT��{j,x�`���Ǔ���(����e�|{���#���i�@�?,P�M��?���B�?���8a���<�Q<il�̣ř��ל&a�6��aRwm͠{��wܥ=��P���p�?׎���b��gcFV��Ňb�S�5�Ap�3��W���㜈�QiMQ�`�T�sZ��/(Lǔ`�����\�bh���u����10n�?q�Ĕ-����-)�lwK��ˠ�w9F��V�vI����_#��,SO���De������|v���3��X5��ټZ�f�1\D@����ײ;�����>��i�ߘ	L�<����x���	���]�z�H��	u�A\F=C��;�:���zx�	9C��x#����sr'p������R�a�j�L"��[U!ZS��+l��/������>�7j0�P�+��Fn\�G�QW	Osq��NaQ��\�����u>�-\�}-J��Y%�:}�����1���Ԙhce�D�msc��Ɠ �U+`�|����W#�
Pm�lg�I�`+ߚy�K폆~��:^q�E�	��S�̩�v�a�X̀�īK�W�S^K��/�\���vC���)�Vq�D�-^ͫ|�zb�ZVDA��q5�x� h)0�,�.+Y,Yz��>����ע;-}"��/�9��o����H|���n�U%���7q���K�l�x�A7�'.q���`m��=#�-�y����sz)� �D�w�}�]wh�$�V�s�o~cgw�y49�ߢ~��y�m��L��!B�r�(j����j������ �m�ov �i��<\����B���w����5�xV�q��X^�$��&�z�X�1�Y�I����0&�Ŧ��Yf�_��Y弞3�,"Ye�R�N�.Q��w'z����Bp��n%r��Jܕ���az�W�Ne�e�T�	k���e�/��Z�++�8�%��-��4�b3����C��?ĉf�.Yh����Ø�in^�H7��θ�	��=V��x�T�;dޙ�V���δ��`~�r�ˬ���q�͏��:�Q���6���q�P03Uhl�x6�䴫k��o�q@΁�2}�@���J� b���k,�ӧA�L�%^+�N���%��i���O���� �W9����*��[�����-�E�t��4�<��W\j�2�"�&�̓Q^CBTqy� ��4j>	qd�9h,��q8���
�E�}��Ko�oE��a�m������� �ۙ:����_Ͼ?��l!��-q�{��m%����R�����Gp`�|����}J`�Y���Ɋ��Q�aF�6��qM�������cw��2��ye�fD�%~nu��� ���Wܙ]��4!{��LՕ���8U�����ә�i�aD~o��`����i+��"ZA��w����'oQ�״Ix�SX�)���'�Z�	-���=o�S�nY�j)bC���(	�=9Eϐ,�J��U�������Ub@��f!?�|��;5�g;dml�qz����s����������!o�	���ژ[�$7ѕ����0����d��0tB&K�V�P�=�$ �VB�����YU�g1u�e?Ysw#����0ܯ����t�i�r��
^����OiL�ʅ7Y���D�� :��=G.�z�ۻ�{�:���;��ā�_�\,(�����Y`G>������w�7y�Ԧ�h꠰��y�ڡ$�g�bh�fy ��i�DO��0�ɓn�1:�����{�*�ɕU��K���r���߲zoi�Q�t�<8�<�=�����	�2:�ޥ)��O)8^(�k�p��av34����̛����2�9�����ֽyg��f���#d�w?o�v\'`�J0���mH�0#W8�目1�4��A��_Pd������I�v�WZ ����Ҿ���,���|��hL�s�o���5'�]�����w�#�<��^�%��x�T-Ҏ��+i=7�"��0#l�q�|(�D<��I�ƣ�ikna�xm�W�ӽ���*;F��Zi׳�>k��%.�{�K�Ha��iBe���X����Ӧy]!�v����r��\r�E\@{�R�T2j& r.
�%aur���m�$����-��μ��G���}�6�M�P�[��B���q2�|��O:�/'��#�1T�w�� �x9��6��:>�x��L�%�X����\|x���vd���X��)M1����m�z�G��VD��P�Ho����ED�99蜢����.-��!��w��,�	�R9*��T���dZ��Q��� c�c0��޼g#kRP�oDL�I:8�����wʍ>�n�?���:CEd��11H=��:�v�,R�����\6���<����b:�؈��T���pjhD0q�!���$؝=X��5d؟�滤	}2�?LKM�-��b���&ƞ��Uǝm�yBsRH��ȃ�H�i�|���#�;�����7(�0�y��T^s�?��>6����B�X	�&�Iy�5nY�@��1@�H�r	���L�:1�^6YS�C�q�`�0�ϖ��4�Z�����QM�y].�����c��-�����R�Tl��{Oˌ6XJck�r���E�N�k4� ���q̉��M�l�(%r��g��QJa�����+���o*�p�:�F�;Qp� xL�T��w��RB@�* ��nE���[���#D�"h��*�	���2���Rys�R�0�Qs��܍ �h��*{��`v
!�e#�CMPI�謅!(;4\S�C`��{o��lK�j8���#ZŬ��@�K��@R��)�B�&�S�bK��R���:$���?C2'�W�\�^/.Ъ����A�7����9��g�C�y 6�:���V
k�d�a�Ĵ�s��Q���i'��;н�ٜ=�G\7����0`��y��?Jx����xBɡڨq�K��9F��Ă�����.�6�K����ڰ'P%U�Pgx�q����^�*NMz�ٳ�\��U��BPv=��y�G��J�s]AO[G���k]SF�����W�m���2\�U�a�����;��_q{�/���R,hb`�vGM=���}ߔ���l�G}�d����u�\�GQ��
˩�ש-��)�P�I��MαM�)"O4o���G��u)�����[��u���R��|+�t��h��Ao��"x���Ԩ�r��Z�rY�����͌�r���`;>���٭``r�$��F*�!KI ܆�1z�S\Ft&���W�2"�r��{�����<�- [�E��S�tk��T	V�@zʌf�@�(��Z���o�耶�NO*h����N��U'��K0/�F��7Y����K�S>_��	��;E}p	���>�ޖtT�$
/6\�>䩳��S�s�U�R,v?�r.N��|��I��4:�q��ӏ�C��>j��VS3�s咷�|�Y��y��k�x�Z!U.�8�X��u|Ab�]~v����B1�NO`O�.]�ɩa���b;/��ś�o�	
�����[$;Z�E��Y��պ�'�Hy�Ƙ�yC��E��'���?Y���R?/�.�F/㋦MT%��y_�v�ęz
�q9{A����ǭ9,�;1l�c�����<ä�g+����0x���^ae����f!q�,K��H2u.���)����U�q��~�;�ȓjC�C�C!�50;I�I|)ls�pܜ��Ƽ^ef����q�q��.U��/p��u��5&�N��s�j��C�α���r@&��� �@QBv'�(���c�Cy���sP�#��=�/-d�A\��/:��H�ۨ�.�^����w�������|`�A���&	s�&Y�����M=�����# ,dP��$Juɡ��ҩ�y:�AT��	V�f�
��U�8�@a�VHg�k?kf�еOh�7����<9%x���vz�X[F��r�m�:��/���PB��&Nb��n�ԭ2K|�p�o���"�	soB�� k�w"�.�R��|��ҷ�JT7YCQ���bw�8*��U{w���{�y*}��/�G�VX�ˠ }�V�,"���c
��ML�%���8G ��D��S���$�J4^YɶBI���o��2=���Ya���~K�bS�h���-J�U:�K8��YrEC^�3�`꘲��2_�a��f��t�t�l8�<ʄ�v�{=6�-�v�+uk駖]�%Ob@����?^���A*�%������@��m�a#*���5쇿�?��̩��vǹ5��͜W�ʎ"RٕG�j�],�0x�Y�����7�Ǣ��'���2ц������݅ a6�� ��eݲ��Sk�q�?܃\;�c�un�_|�aKxx�7���(|�4��jk�w@�n�o���I�HZ��%�{:�J�hQ*#��a��j����MW���K�-�4�I�Ϲ]�|�����B�����N=����)޳��LW�`�"��G�b����u���QN���}IE�TZ����%��|�� -��<u�j����1?[�T��ݮ]>e��K�㫞�a�WS�p���x�X���X���x�(,El�
� ���I����H�"���\�?;?Ю��cE�e�`[�W�??mFJ�|k���#q��#��o��h'���W �4|D�u	EJs<9o�������*��s��UHKs j�硁��7�('������oe��_7�ic�}H.8���M�{�_w^�94_�hv0(�Ju�k��I&���c=V��ND�# u�!�#���,�,��r�;�F���7|��{����NC�G�x'm�ui:�Z�Q�� `����[��]���Ue��4��Q����~�<�V�r����T��1��U2ԯ���E-Z�;?��1�
�Δ6��J�����g�?n�;����u���kg��5�z�Oy�흹����f���w�ıSY��rj���?Ҽ�v#R�M-�$|� ���@h=hĹ�+�K,��4i������G��$�X��a�5�K�,಍&<j�oȰx��
��R�i\�r�y�~;Xr��#:E�	J��D��v�Q&"��1�}�����ӏ�r�:�@D��0�1J�d����lR�R��ΐ�������5T��� ��1s�g��̔��h8~҂KFX�Kv�hK5/:��|t<���ǀ�.e�1V�=�ah4z��>�ՆnO���f(�OW�c�C&�d��6 Ӥ��_�a�Q�/2�_ܖXa��u2P�;�`�d�[�����q���>��k^�Zop���%`��� �IF�`�@"��i��kQ�Z�`���mI�n����ku�ª��	`�ѯƮ����¢R/+c��\�V��&[��S%���n�^H�;��V�b�<K����~85xRi����ԱB!B�5��e�r�
�ETe%�l*�Y�F�ၶ�~�^�ц��~�G��}��G�%��F�v��s�������4#���tx�m�Ϋ���2ѽHޖ��)����M��y�S���=�������X	֍^W�Y�	r�c�.���tx��K�ASX�����	_��?��<B�,����@����ч�iD��"�>�����3 ��+�o������*r����<�ߥ;�(�~v�`����#��6�J��6�2Ԇ�DǪ���ȇؖ ���#g<J�����^oU$�j$N��L�����k���y� >��R�C��i6�ɇg;�h3|�6-���~n�Cu�I�Y;x���E<ъ"����]���!�,�PB���#j�Ӗ�fn��"�HP�&�#�eg��>;}m��~߹;���:��c�.չ�*C%�����m<�}]�,���w����8�� ,N�KM��XT����dq���"� z�[W� �Oל��@����d�T�s� ,B�|�����X���twhW=	��@��M���;);�:j�8S�ٯ��؃/OR�L�����+�;����D�n:Ӎ��BE�k~��5�rB��J\�I5"J9���j�P��"ؽs
G@��ra%�q�}{}1}ih�9�����!������7�2�!��o�6/��O��s[���9YB�;��B~�p
2�z갘�Y�1��8G�w�BR��b��R�o~�*�y���'���!%&e�RHX7sL`h��Z��v��7a���e���̮t�"M�b\a��r�m~6omGT�6/X�Ӟ��7����(#�g㏈�ڪ����#C�t$�v(���<p�M\���˖+`�Ê����+�0?�;���Z�Wٜ��G��5<��S�e���m���'lڟb#���!�i�#�_B���+V<Ӛ �iGk�f"sM*֏,i�V @�yU�,i��<-�6���>叫��j�bFtPV�~285C�Y������A�|�g�v��R�?��?����\Na�+��F���~�3�bX�Se�Y�xy���H�Z�:c>0�F���So�6��L`r�ϡ��$�9qrRN(�W��{�/}�Xk�5�(��:s��|��%��y1M��$72NiF i,��>�L���+�J�L��θ`�;��E�63�t/�7G8����װ��o�9U#�U�۳Z[*د� �6��?!n�-���/;��^���e��:��U.E5��C?����*R��Kǲ�ą}CyCpTҭ �8��o�Y���������mWK�f�������i�>N��Ȧ�u�}��~n%W�4��Ā�n&�,޶-,;�#Nz�X4�Mf��ǚM^�ӑ}�Ȃ�-BG��7�R{+��᳙�]�
�|{{� �v��p��]��)i��%��<����Ax�$�\<�7�����s��>[�y紩t_����S(\
�3F��1�ʅ��� Fn��E988!i�WB?!Nۋg����蒍$&X�i��8?  ��jCtn>mvws�^��ω�t��S��P��N�'
EOB�^����܎ټ\Z�oJ�L�jEi��`���H@�a�����m� %�Em|ID��3��Q�LaZM�DM�
�@`�1�C�kۻ
�X�3	�������`0hFS�mμeb�ч�B^z�``�s��pB�J��ۥ�2��y��Q(��Z����R���a�tS�);:pe�a�֠�ס�A�6�6�:X��������K�%�c�q�\���d��6�rĦ�C�tF�R�%����\�X�m�\�-��ɘ)����}�@���evch�$������v���;?�W.�Gt׭��g�L����������X���:�����*>ًH�,Ue:	����/�m:��970����Q�T���ׅt> �ؤG)�P"��:�go������U�sU%;��8k}k��P�ZW�Q�ɧq��k���oy�ķ~��`�X�-k�}U�B�}�������¶�⟆��p=*�>�	��\�6 =3���p���&o]�{�s���Iʐ��=����[��Z�:l����Pی�X��!)��=v0iኧ�* �3�8��8��̾�ep�g�Wn��ڶ{��~۸a�%<t�#x����j���
�g1�d�������S�E@����x��z�_M��_�	q�*kIͧ �V��ΈL
��!��Jp���x�ՠ��CvZ��u��xP3y_1�֠���J��&~�*�0���q��1qr볙���Ύ��+�}�u!�7`0_x|i����iA�z
�U��$���R��͵����ᣞ܈9*��x>JB�l���OW��c�� ���!P�4]���۱#�Bc�C���c����Ώ��:vR5��@xtv�V݊G5�O�;��$jn,9~$]�wmЇ�lAPC�:n�ׂjA�^ m o������D��F`(J�vk[�懓A��nuq��}����� μYO��qΎ�h'
���F�u��l��g'��n�E��[��t���j)=���=f!2��?���)y�rR�ƦXQi{�T=�D��`L�X+	�N��:$�%��h�M���J±���"Q������pPb1� M�&wJ�$B�u/a���hM"!5z�a4��:�Q�H��~�W�آ��p%'UH�]P!&�%	�ZF��#���/�	�w���t�9���gu*�c=}K?b��>��IL
�%p�PY�ه���:+�U��S����f{�+E;^��)�g#hٷ�քwI��j�Y?�O	��u�W��c,�t-j�^����b6�˯�l��x�9�[e�_�%)-�ݱ�Y�v����xN_�D�J��#���-��~5;�շ���L~�Ms��6Ρ�<���Y7��
��Rl��� �t>�j��`�\e��a�q�P�#�mf��H�D�[fآ,H��4��� E������Ə/�^����M\75�<g�,�%��	%������?����癙$�8�4f���2
,R��m��	6Co�w!\(5H5*,��9���Y�0���wme��B��('-�q�M�J礱��8U�W��� ;�)4b�T�d@��8��T�ȋ���FƏ�ӐY�C��a�)�<�"���hGD�3R�z���`��z�=Ev���׾č��sr4XlaV#��,]j��{B�\�G��U?�'�F:n�m����{��jD0�������{�e�j��5R�0�����--���Ňϥ��-�E6ק�}���P樍��u+鳐�'�Yc��9^\lj_�T*Rc�P�6K3Fn�ꅼ��q,µ��8 3���]l^����<�wr��ᰖ�넨ef����0��T=.�f�)�{L�ٶ����~,_G�9Gc6�Oۙ{J�u ����fK \�%�F���g��>�֞{�F;���(�������<v�*��0����3�uY*T�J��%L�F�qY���^�4�.5�]��jx�@ֽ��#�#�\8�����#�E$f������R��ߠ:��F/�T�|/�,�B�W��:�R�A��V$=��MY��-��|�f�y�Q`�<[n��e��o����MtM�'.�QJ/�&={��C�N::�a^X 3~��=n�@�!� �8��M�� ���𼧹�S��b�L���z�0��S�դ3��2�" T����1���#�%�<��1�K�2 ���2J�]�R��oV��%:�d}��$��*��hq�H��;u\�q�	z�֕c,X)��L���S�T�i�+� Pݓ!�� _j�����-�r�3�L�,�����z���J��p��9�M�s���̆ .�V<�){sb!�]���]��);�=��� k����W�<����i�أ����CACY}�Y>�d�U�χ����F$��p^�FS��ŕ�klv� H��U��K��g����m�N�c�a��bUu̹tޕ��-xGL�5�0�<�Q�{��{W�D���1����1^Ea��f��%O��I�>%��/���#aO9�}fy�Z8S����H�4���O���^��p�K����CE]>q�*�#p6Rq���Mَ�����ʚ��\�O���e��"h�-�T��X��H~����s���'�b�bK3ِr��C�!]��ڠ��O�=��m�~>�+S��q ;E\�����e�i?y.!�2} i�Ѥߓ��̞����@휢N�[�Mup�_NK`91(��n��0��7uю-vdԜlp��H_7�a�������G��m�TY��@-8)lN��K��\;ȯ�%��Nk
,9�%�wIn�g)�-����L�r�!pl���3��;���j�E�E�!:%FW��D���R̆��y"�	��4��ă6T���=������l�YZ���/��c@��+r���V�K�@�]�HHK���{9�N-׀s��>������*~$.���!�ho���|�aKz��L?m/W�P�
�F~�JjG��N}��ќ�40�۫B�e��N��-��8�t,�ݖs�=�+Zh��xA)�}M�z
f�>2�Sց�-���Be8�z�*�KQ���+��(�stG�|ؽ0`G�Y��"�rT����[�@;�sV���	���c���*��x�t���6�=}�<N�����2�"��|J%���[�r^���Q�Y�ci.2��Uu�� <�Ƒe�g~/]^��G�Uқ���U�/2��'�QOz����H��6J{a���"��8����Hm�u�(5}v=����MvDW����Wk��~hl�� �E���Z�0����B@uCs�_<s�o0$�rNj���S�d����廓<���R-{jn�/'�84T:�Ğ.���̹��m�|N��^4�9#ɬ�RD3�tr�� E0���g���3�'f�6C�6Mg�P��Ӽ^y&�ˁm�˂ۖ��`��̮��	>��̘�'�[�`QO��j�A_?�Iv��u]Ӡ�l���%E��2�$�X�ŏ���d��;٨F�\�Ĭ����*k�a������K0ƹ�P����%w���h��i�9S�L�g����<Qx��^�un'H0�����{�	N��cm�x�V�R�7f�D
�YV2���!����g��X)".�@��������`}��/K��=��t��ӡ�B�s��z�0��\*�ax�6�#_�q�^Щ?���L	�fj�����|d��	Rԭ�|�蜢]�;2��������m��]�_/��"��C��-��S,���I>5�7]����*N�+�����Ƶ�^b���46��z���/���)�+�(S�:/o|fۺ��K�� �ZH�~�ͰOX-����K���iƱ%�˂�@���`�}Q#���P/
��i8H�{�\�t'�Z�1/%�˜�*u��O叴�^٠E)��|��iy�Rvk�B��(=>����t?��w��\n8�D���F,v��ߢ>0���m�*I��'��2�D'�żմ�٥���'�DşIK6Hl��x�q-��5(E�F>�P-�
f����q��A���x&�V%W���'ǂ]԰��=�}E��>��X���XW� |�a�3�a��o��Zh�6'����y�{�np���j`�M���I�V*��{��ƛ���][0tp�`gs��
j7��P�e����x�_����D ^/|ָ��)_;6�*�W-k[��Mг�u1�Ag�f�s�P���p8.��zZ��9��[.F�͞��R�'���6$>�*���k�-��'���< -f�U�}?2l��t���n�h��^�]�J#�,^ϟί�K������ϙ��8J  �f�[�NJ�`�%�c hs�g�Zl�$�� �2���g��	N19Q��ݹ����G�b��Y�^���Nn���8�,x:^*lsE��4
�DTp�{x�y#��|�]�^���������q����r��Dt&zw���,��)���g[��RG*��i�f<q>��L�0O��R�_x��I���F���e��&�����P�;H�jϜ}�'BU�/��H�Q#_-ϵmC���^�c52�;d0dj�#����Fb�]�w�M��,��69������]U�k�׉w�	E���۸bx�-���TW����/�<�h�ݐ.i��� ����ȝ�Z����m��·!GO����4��s�o�>V�GQ* �j�i�Iv�qܷ8�h�8�Q��~ŋl�=w�}I�<Ȏ�!z�C�6@�t�2�v�����&FA!݆��J5�����^ ������HxLgA�������8l�UI@ά�@S�^���u����7u��W{�#*/m��y�y��e�i�o�]�]8�����-�8w!˥@��
;���=��ˊw���E�t�k�b���E�pEV�T����0ּ�<�2����R^^ �G��8�1�\YX�����T�w�ޱ��,�x1f�F̑Qk���g��C��6t�>��h�-܉̲��@�2�؜'�a��:`$n�TXgY[�������*~�T$��ठ�_��w�'��a�<������y�~($o��6�5��i��0�p��H?1��e$�iQ	���c*:�~��j[��_c.C�٩g#���Ѿ����T��YJy�a��+�Y�pg ��ǁ��h����}�ir�� 6Lq7�4�\e��e���z `��@��"9��ʭ:�K|&�,��JĊ�]����NX̖�zJ'�];����3�h�:x��G
�Z���tX(�8���u�.~ݕFst��v�p�a�5-c@�y�s[,�*���k��(G��ڋh
̓4��m�٧w�B̴��ن%����2�d�r�tc�˸��^���j��,��?gA ���/�k�a*�S�$%����,&���j�W�o��b�y�@��aC[�̒0i%��~E���e|��aj��"��:q�n)��9�G<E��rў d����y��-T/�_趾�?�QF3
j��"#�:���Vw&}��e����"��������HJ?H᫵Cb<�ng���-�szP[t<�1�vT�0�L���D}����l_��L���2I^zz+����x3=�o�kIڦ�$���B��k�2!��X�+�M�q<���K�ա�*(X�&v{�������ՑC�Q���TOA!��hN�D�����ESV������߉��� ��6������ z�Y����sT7���t%ݮ�庿F;�gT�&�7�(%I1N'�K�+|��G(�"�߶s�+����:��Ќ\c����9H��*�M�Z�s�1��|'��}��|KE���bPpE���� ���1N������=�5?�K��C�E��&������-�|�У��a$�����B^̩ѿiI���@N�-�,���.��`#b&�.��*5��;����
4�ۤ���-Q7�1�� ���Ӎ�����E
�Ģ�Ħ��He5�X5e,zJ�ϸ�J9����x#a�ߙ��P����[���I,���S�3��Y�I#�(��ϻ��4��9�F1iw���(�B(`�� M�}��dzp��&>RE�8���h�ɬ�S�=�UwI�YPq�[��
|'��r^�o܄!m��o�#�e�Se{B�TJh
������m���&��8�s��ߙ��	��:r�ra��BU)�ؒk��N�����a�DH��!�W�3�v�aa눃-/%��)���1Eҍ�]���'L�����\R��px`L}�u(a���;A�|�f_�=�v�f1���|0D�����yS��y4�s���^_�=5$�瘛�*����������]�P,�<ۙ�DJ�u-���MO^Rns�:6I�C����[�E���Q��į�	U���l^�4 Jɦ]
��[W�[� br�qk���@��X�ީ�����v��壄v��C�$��K6�;e9�A�v�a�j.�5���s�-�:4��^2R��eN��>Æ=����uV�ގ�DWF�8��?A��hTla�v����.Y��)�d'oR�$�K�Bގf���F�+�F�V���:ޔ[c��~k��tG�P��Ic?;v�����~
�][�>����mL8��6x����6^�T�Ý3�� K}���a�p�'yK�Qf����1�"�3�Gz�J%c��NZaee��no����q|ξ��[<E'׎Gz �J̙~T��K����Wj nN�b��H�|�8�|�|��z=�KQt��hط�bs2)�d��D��E�^o�70����xo(���#�D��ꌱqU@>���"L>l; ! �H��>BX�0�o��Q��䎬��A�� `o�n�Pɶw4�?�L��e��hr[�S��Z�O����E�����1q�Ni:��)����t¶�2%m���D����%?�.��F:�S�5w2n�L�lZc��PW��",]�BN�G<���4�ˏ��Xីo5l�����<s�5y�l�+r?ܐ���S�ft	D�B�_H"���v��,5�����w�s��dG�9�� htΤ3�n����D��#�O�5|�XO@�S�P4:����!��@o�M}w)Z�ͼN� ~��.�Y�+h%��|ł�c3��W��xW2�YKeqD-p�0f�Ks�'2��4�L3beֆ̑���r��^�S��']����~%S�N`ܚӿ!e������NQ�>��'�s���x�?�5M����:�m�}�fX�+Y�MH�^��,�\^A��&(d^����nJ�=E���D)
yٜ�,B^�yy��u��
�L�ɵxn��7��5�2�F���hs�ڴ�&�	ڰy����l�(qD���l��"b
�G�%gA=׭(��dE��M�(�@�fș�W�h5�*=Q�h����Ht7�^X�8��r$��[�)�;���˦w(@��3���6s�2?G�(i�&q�U����<}�	C�F��T_�$ƀ� ���Sr �@uɣ~A���0�<g��˻1!M��W&��W]��dk&)�5z�:C/��p){�m��;��wB�����9V���Yf$�w��U�
>^VՖa�;��gkCb��RЇ�'�ճ�f$J�^��L�!��%�[|N�'�W.�I���@�C�d,2_�֠)Be�8V}����'J8L��כ+��gjx�ɦ���K����*? 5,XB8N��p���rk/*u��R��U�|TE��L�oHN����Ļ�P�8������ݑKF���+�����z�b�������!�3�����0����#�)2�x���!)��W���}o`�\V/u���N�Ni�c8ed(v�p�dJ�����{:9P��$$��F��`x�s}�����]il��� ��T���h�kp��R�f��ZJ��ɘ�X+8��vi��$�
�����II���� �>����m��{��c���{���48�R������2����X ?`�9��c�/�[����r��y;�J��/�l�C�ße�f*h�d6�de8�!4%��Z��W�)8ըu-A��c��&�x�������T��u,b�י�U>�t�)Ç�C%k&��/�	��� GP)�|��P��S&2~BT�2@���z��T_YP��$,�]#7��i'>3E� �2����A~�9�j��r� ?3�/C?�O ���U��P�F��U���Q<b�E��vi�ƹN(Vcoی)0~�s�<��MU�E_,�?��"�@Y�E<Q�1J�q�v}w�t�q�����繊Kn��{͓~��?UXh|L#k�5@<�����]�ta���㿗$Z匫	��H3�c}6�/0�r��B[Ny0^z�h:yS�"g���������a\t��+a��~`^~[t�fb�R=��j@�+�6�m$똱	���a��f�x�U/�}�ОK�!e��[7��X�z�u��{��f�)_y���E��Q}\��w��5.�������?�s���/(���%L�X%k�C��n����4�e����7o�/u?���� H_h����U�@|d�%���Y�I�нג�n c�g+����իu:.��9��!ԩ ��Z�����C��c��MM�Ct��$,\e����zp&�]67�_�����X�����i��u	3}�߇�����6��m��$G�*l�z>R�H���L�/���Ӎ��S���p�"��$���w����Q�l��9����B��-�o��9\@2���'`1���s>�%UIWd��ݻF?˚��E�yJc�-8���5?����ċ�ѢL(i��Q,��D����Յ<�� 6e��Ap:�MM�}�~�gD͑7�U)�1CD�ɨ�E�����\�"�%[Ku��:r��}��^���%��*-)�<~�P��{UX!�-�&ð�k��Ri�f��O[���:%Sa��8����R27��v���5 �_��ރ/=Β캎莶�X���r]�ӗLCc�tr���,1o5�Y�Hm(�5�%�j��@o��n�Űܗ�^��iX�4��`�#����&�@c'��>֎����U뢐 "��>�ˢ%.^;�i����le�"�����Pqip�G*jP�� �T���)��O��qYg�[	��%D<^O)�R�Q����P!kT4,�,��[M��`��.��:}��H9*~n���6����_����p�vyg��F�����Y1���t������Ŗ?����N��)6r\GU\"����`�5��q1j'��lyaOly�����;�i�M��ևHrxj�W ;̡ʎ5�#uXg���~Y�B�G4֤}Z�Y��3ЃS7kf7�9W>Z��v��$?���榇��a�<w�$��M�{�9�kl&}��.���f��Rx<�����+�E�"����@��ͭ�zK�Y������LeƉ�X�P�
�ڈ=>q2el@�o1I=~X�P��6�c]�{P���خDM��W\iz��ƨi�p�]$��f�vP��@�^�a�\�S�##����w�*O�7�����L_Fg:�j�J~L9��-�b��{��&�S��6�.����6�ָ�r�Z��do�qï<��|k�c�i,M]#���ڟ��������(/As���S<3����SLr:m&�qvrk9�4�vS{�iI�蹓Dۼ3��j�7�,�y5�^���wͳ�F֫%��ip�h^�*gW�؄�/d�s5׍��NA�W/�%;�ۚ9{y�?'�z��tC�����z����.�4JI<����MTb=["dZLpֽJ�q�=��h�YBϊK��v/��W�H[�^]4�vɜ� ����&� P���P�{:����y#4�b2�[5�Ӵ���9�`�����ؐT���f�X�_�X
sEֺ;��+ &?N�P�$?����f����Q�dln���o��eo��d0W���g��.k,�5�����HN&���ڦ(޵�i�|.6����XG�� �R�ϋ�QJ[.�8.'i�ksn5�ȯuX�~aB�b;UM8���̏Ǡ6�h��!(s~#�W;�+6bN����D�0k� Q"�<A��=p�GD�'�]�'���O|	8`��*�`6v$=ke^�L�PC��j~_��Ư:1�W #}B�d!��us�t���������Dh�5 >�=Su���PǪ��7���G�b��MR������<1���匝�y�COe���c�S��Ŵ��j0£�A�JN�j՚��\�ǽE�C-�-7l3��S8B	Y,f���2��kL�/a�������/.L�mg�t!`f����*ڔ�X;�uFm����QB ;�#��DD-�'�P�v	��wz�ID�B�+ߔq��5ʠc���"�x����%F����*��K�3�(O]	��a: �s(83
���M�pON%*d��#ys��{[0q�7=��b��E��G)<�ٻ' �*x3�#z�����s6�pQ�|'�wT�SpH4��&͐�RN5#��~�)���G�q��9iM�+�~�j��FZ�<
�������"S�d�KlhH���=�FWN��T��U�Q�nCfP�,�.u�.>0�[�%Rc�m~�
�QE��:�����ҕS1ѫn]0|���ѳ��	Hxf&�I�� w�mF�������%��z��|W�v�F��Z�+z���y��pA���@*��2��,WٲÄ��a�V��!-L�f���
UN�ʍ��ѹ���An��T�-�55]!S?7��l��N��O��w�v��ۗ�U��0L~�%D�!��r����ܮ"XC�L���۶!mS����g��h�~hz!�7:�v�-|�=;�&\k�e-2�3
S�p^��!�/�=*�&��g��B�������9{q����S{F_jEB%�쪴ż�9kHu��BOH�\ذ(d�j5p�)���jH�'�!�D��
��ܾ/�i��7�� �l�.P��b�5�
cqN'^��.��2f��Z���q.�&�J0�j����32 QьC@\�=̭a���)+��yn�%Ƹ�����Q�Z,�� �Dܖ6!��}[`�s�����MK]�*����2f��|Vچb*��\��8����`=��;Bf��- 3�E�>D��֯��$L�=y�was�����-��ط�Bnnh�p�IÒ�t�����Y	�ϥ eX
����Q�H;���ڷ��t�jpo�˙n)6ny
�gE,`(�>K��|�_>L�������0%v�B�#6z��J7e�.�RX`k_�5Y��	���^�sA���5DZ���JH��s��o�y��3/��uwo�0Rn�@��-kI�����A�9c�z��2,r�@V�1�ZOK�(��Z
~�J�>�}��Ȟ'$��{S�����?0�G);Qp�°G�w57b<���Z�Nz��w�ii�*���	[2�&x�a0C,
 �>],(�hx�p�3����	�p���X��&��V�*�*�{2��)��&��p���3%fCz``-w_+f��p*��gR-�v���?B�f6rJ-��'o߷NR�^���zo�!h��1;k�tc�.�H�hh��K��`?�(z�����JӭI�Y!�cL>�p*2����p�)z��S˕�;�!�ʊ���}ܘ �2�.㥦ľ�B�Ļ�F�M:��}IGI�o����Oɡ�dy��B�I�̶��5 ���cD��$�������@= u��(��X��e���$����p�p�^�߆��!����S�-�ժ]+S1�B���!y����Z,�����K:;�]�㤛/S�vKX�q�S#��{c�^6��,M�7t>��a���@���� ��'�##��{��+�D%��c#�^ (��#�+��}���؛��g�k8���L�Ǿ̇/�R9Ԅ�=��~�݁���P/���7oze�b��M�gq�@��;MR:��%m�y�{�ً	�5p�8Q��/��3�r��������.���,;���{�'�Ү7�N���sV��P�m����EC�T"A�z�?^ث7c���Mm��i����NC)�G���::}$����7WO�[C��v�h���ۈJ��D�RA+hh�9Z>�18��y3�{+d��:,.�pZ��D~ �b>up�b"!N��<s��d>�i���!�>�и����>h����P�p�J�����R!��	�|qދ��i��4�]�Q������BV�}c��&$�qJ�Q��W �D�;=��W{]�BG�6q��R�F\ ��VE��>�
�'���y4��V:�o�+���]@i�*�2|���M
,J�Z(\��!%,jE��H��;]z�<:n�\�C���h-ݚk׵�%�r�m%m8�F�"xM��iH�e�<}T�W4�aՏˌ�Î}?�Qe�����5�̯��A��L�z#X�[����sn���>՚jU�H�E��&.��|��p���&��#c��_@���O��O]h�¹\Ɩ�jn��]�a/МWr^�йźl�q��K y�����R����h�۷�m��'BD�>�ImمR� �-
�[5��S��,S׮w��	Q�O��WE�B&R�D?���c�����'��z1T�/2Ɇ� �;�_e�L�c�̕m���D|���t�/\�{�l�97=֋GU�A>�0��ṱm!�T%b@I��������K\>�%zr:X��]�E���\%�(\���{��E�����bs3��m�7��h�L�ꃧ��B6 Z[�_���5��8>�Ӽ�OwWqC�O��rZ�Xu>AN[U1W �H��0�t)_&2�Z�ȸxŁ��r�o_?v�/�Pa9"�Dy�G��U��O}�v_�O��i�Ѭ=q�����h��
ORF��>��s�X����������$ۏ5�cђ�s�@�3YXp�N� ��\��� ]��oVG����ى�HB�e���t�l�lS$��B����Q�U��g4�GVt�M��������6�h&ji�V�h��]*~vZ/�
�_�K�H*iָ��<w"�&�/��`;���T��_a���I� &BK�Wv$�75�H�`�i庀ާ_��޿fF�]�����u��1-�@�+/m,�8��xs:��u��3D]u�j#�
������f�f�̀�H:�%g��j���*�]�iL�y��ٝ���,b/�8f~g��(aѫ��裌FT����Ϥ�q���'-�UL���o��\Z�6�u���
	��+�y�E�r���b��l~�vSq38�C[����LzA��P�ї찭C<a�r�$@�$�t���"+7A�J���{��C�>L�m7��5|6�S܁��΅�a�N�ߖ
;�h���U�xMi�A��&eNFw?���	����ޭ��ᬒ| �5�ṻ �$��|���/{��/��DaY&�
V�y��NeE5oI8b(��~1�wiz�e"v�a�_�J�눢�!����X�������0o�#�+��-M�v�.��/�
sGϛR4�E�*5fA��C�K������o�_���Sj��?1�q��6goa��K�
��u�W�@5�ژ���|<�X�S��.������N�7>o����	qQAT��c��Ů��D���㼙v�_�Vo�ͯ�q.^"��۬��8�<j׽�%z.� }��~���#��Wk��qL���m���2����sA�>��`�6UU+E��}�r��H�������Qب�+�(�5dq���2	��T���#'|�w>1V��S���HI�F�J�~1U!�>�0��$W6T����I�c�+G��\�c����%ܻ���~��x'
�/c���d�2��9��fSO1�H��?Ĝ=g�t;U91p���_y�ށB"`FEP�	W2q3cI(93��RR�w�p��k��dӓ���Oe7{/�P��hk�b2YU���*w�V�ѭ(^��^�V¦�LN`�z��o�BʇN���B_JƢCX^T��F����c�z*_���]������S���%Ke�ǝ�r���_#�g�vY�`����mtz\̴]�㺦��y��<�
�V˯�a �:�����mcw̧K�[pz���'�Y�rF`���.飱�c'�ݕ�����`�:�5��5��\�4\��Be{�4'=#/���=T��Y�^V�X�g�76�/	��y��<�*<��Ԡ�ů�	�qya�9�}ڔ'���]���\�c��Q���XA�/���0��tK�`�UV�ݥw�pO���s\R�un�g<��4��u�`�������	�
%?�@=�?ج�?+�bM_���*ʗGph�Vp��h�6Z������ʼf�<6�=��7�M�M��c�[%F,ҥ>�I�b���BrUC�@X�c�q��C���)�v��+J���Ӯ��{�Z�*9?�I:vF"{qӲg�T��(ְ�d���f,з�b�x �w��SVu>��S��ӫ蹷��X������ԭ0]���\B��k�T��oƖeld/:����1�⇕�%0c9M�o��N�1Yn)y�5I�e�F48�M)���v?�
ͯG�Z:�������e�9Q�4���3������rvv���T�|W�x zUA*a2��䎽�#���+N��^/\���w)_m�hKr�}F�fe�YI�H�� �$�c����bo�.�r,����(Qt;Y���3�&���{I�
��D�2�^�u�f�g��;u��n�p[���.sUc�eF�Z�\A�nJ�&�X��:����p�F@P���+��iI��-Oh	zo���?J�V�!E'��â�VC��N��7��a��:�{j%�X�q!!�
mFQw8����=�����#w7�Ø��3d2���#&{�A��<��u/-�Epi*�+!���8�#dN���U"�2�$�
�ů���J�OJ	ǁ�*0���3blK�evAm��l�䔜n@���
�a�-�e�;.EDF*�KS��]	C:��(7þ6!Ӈ.���)�Y���Pݙ�<-�]n�I
Z7M�s�-���vkʇQ&k����^����I�o`P�Z"«chz�Og]��c�W�!�{�l�~e��e���b[;u�Ծ��M&���l �m^�'H����:�@H���V�@�,��r(=���x�mx��Y΍�8d�#�4�<N���@s�n�����鐀�h��])K6�ے5@����t��2н't��h%��6��x�L�V_h�Z߲�1�@	mh�i6��@���]��1���5��H΂�� ����I=��yc�考y+��h��Dϟ��/jm65I X^Gx>��?�!�߮�4K�^�șyJ�=�B�I�`��`�f��5 ^.F	@`�¨�1sߔǿ���>1���#���\��ѶQ�.7�*��#G{�Ϣ�h��>	$8rQbt-�Y޻���Y�xa����y/u�����{U��3��@ߪ ���N�~�A�5�ZU���t�yX7+�.����0KS������ ���6n��Urŧ3�p;z/8w��U ���F �Ӻ�/<ی��.�u��6��h7�Y�b��� ��/n�z��<;��\�*Vj�f�����2c�6R��kG;7����$��n��Q<�9�����x�3�����	t�(��q�'
5&5�_dU�2�B�$�l�'��Cn�꼕��vtP�!���l��2��D��ׯ1D�2��
J�����G�'��`��u#o�]�\��{E~��-h;��s�U����U(UjQ�1_���{��3'Yt��ۍM�g�g&sZ x�4�/��G��
J�W�0���㥴=���{���eZ��H�:���֖��V�il7�����W��M3̋hd���֝��V@H��W=��rͨ�N�;�%U'�r��W�����U`��L��0� Ɉ��AxۓE�I�pL�ݯP��y���	L����O��������4}p�~�'���Y�A�oZ%��k�YdG/ �.� ����7�j�o׺(B9���d�A�SV=�����'���5	��s��T7�(n#\�����+��h�:~�5��Kڡ��4�����Ҡ$/dQ}��r���{��M�������0�lן�0T�|_:ܡ��fw��z|�?�
%2�#��� 苳���h_E�Q/3U�<��\�%$Tj����r)����w�{��	����7&�> g������fR�uO��,�-����:��F��R�VZ26�M���w�H2Yw�k����̱]��`kCL(��9�k��%�W2E���\ٳ�{YCHC|/�~�sb�~�����6C�n�˔[��p����7�ܒ��}�(�(�tr)���8c}�7��V�G���#nV��ߴ9ޚ $S��DK�ӧ�qM>�VG)DT�!餺�.��n}G�&&�Q����&4�و��*B�i_�:�p�~e9� �����yWM�ߟ��҆T}���
������U2	9��v���}���@.Q!Wpa�{�:�!��Z��ZE�G�l��OzOt��R�����f0���u�j ^�Q��;���.S|� ��+����o[��jS�v惟N�?�����9�Yl�ea��$��qO�@�<n�����r���>�օ�3\�E����J;ϰO���tr��AY���^3s�p���/��wW|{.�YdP�Zi<���\B����
H#5��07���K�w D?�6�N������W�sK����D�Lw�����f{8��<�1i8D
��fwlT�B�|��
��"@N�.!�u\���ba��sё��w˃*.h�]I K6T����~j�<� �����YcD2��&��}�A�}���	��y���Y���ȓ�n�	:cCW}�!>Ea�f�ɢO�4�ͥR�Ѫi���${r�F�Z{�?�~'�	s܆s¥#�{�쐖�������l�A,�p5���e0:z��u�����:E%����1��h��/d�UC� �3�W����Un;l8�)�%�87�����������(f}��e������zT|.�D�Z���(s����S�J��^]`�;ڤtZ7�1�^�
���<��L�̵�����]l�}�J'�ϰ@p§���vg5�Ad�1Sg��T�fH�U���bv�^��T���0���h�]wu�m�-�{' �6ׄ���c4�űܚO�t�! .|�4�OsSG�B�����X�]h���j3z�DB�d\��-2����V��m�+!����X���e���J*
X�����L���/^���_L}kH�e`��Ѹ[m��U-8S@��Z��L��w~L$�xt�a�m�u��>�_W��м?Z�}MgX�6�2"W�rG'�w�3k3[� �O��P/�S���r�ϋ��C�� ���][�op�x��/������{����T��-���v��U�%�d�����aB����a����u���"5��O��!kJ�,��?�=�ɻ���ƌXB�V�g�7��Q%�$K������a��5�U��?�zE��HhKc#�fI����0U�; �⽵J�N��0���t���Կ�M�P��3�@�/�=����f�,�goT�@.�K�wt���㋺B5�J��a�&�Μ�-����O|���&"�t;n�cxZj3Z���9�#���:����Z��ʗ�6ҷ�{÷��� kN:W<��g�
��X-�������M�vNp]Dc}�#͑Bgeӕ&h�6�����q�f<l�i���:Hq�U���)�&n�������W�
�4��m���lkvAJ�9H:<�#ws��:���6T�o�R%�N�Oa q3��q�Y������?.o��� T~.���֤�4���i�o����@Ȋ`p��0n<� �ueJg�T���Ҁ��S�BC�2<��mT�bW�1�Bw�Y�\�8�GhnfO/j�$*��o/��yE9q����ϗhѯ���'��"��r�,N�^�N>aB�O*|/�Z��DZ�8�	��D�#~ȸ��^2G�����xc�&ra ����R�Z}���I��UQ�ZPj� �{��tZ�?.?�A�9*z{ܖ ��Z#���c�AV*+�"�%��GS�Q�ń�������l�?��#�޹Ԟ�:���Yw���!���Cb��?��lT����A��5s�f'm-����)��m��<2��Dy����w>�~�T��Wr��(��L�+�iG�a������9��ynQ{��$��r�����N���?4��}��k�>� 1-��}�J���:�P'J)}<ɴ��B��44>c��x�ny�#4c����/x�s�Zו��|㕠"�,D����)��]�š����c�F�t�]
M����}�܀!�LڢGn $�F^j�@�'ٿ��[��!��T��	�5�7�j�n��9�N�!�`k���w���F�:L���r.�[����h_BkHW�a��2�No�'��Ü�i��Y���k��{MKBw�)�z���JR+�^�0_E5��*�d7�tP��ڴ򆼪+k<[G��G��^e-�g��ǋ;��f#�'�9K�����.+��+�+��I�����m��(G �/�.�g���!Mo����qַ�n�2uT��J�:��	�绤V'�3����G�ٓS�:"���{�v��9� V�f3�\0�\�xi��sLn������̯��.h�R7Wilif��K'~陎�� �!]W�}�Ջ��=� �l<����f���.+��(�(sM�A��y�k�6�S��љA��7�B� e��M�$R3��S�q^j��#��nK�]���6��=�A��� �Op�g9�o�5'�|���=ڀ+c��b	8�\>�m�0���D��t���X�*��	W3!�h%�{W���ό��e�َ����N�\�C0H��s��J�~3]�,����:�R�(�r�@KS��P�>W������5���z[��"�^�T�Z��3I�������K^Ghf��)ʏБE҈#���]۩oX���O:��^%U
W�&��.��GPX�p	�|��y������7�O����w�3节J�I���zW]R��v�Q�> �L�0
�8���?FS�a܀d�X��p�U%�V��#j�Jt?y��_t��1>��޹٘]���M����R:!�@���i�7��"�׻��bD�>��g���<�k瀕��{}="�5]�Y��_K�vw�+�zW)Ab���=W�2�v���q&�ܠk�g50�����X[��G�"p��Y�J�"r�g�t*�Z!$��ն���	�갹����E�.��#��ʡGr_��^S׹^)�GL!2޼�խve#C\Ր9��@�I�hq�Ǔnc0Ǘhq=�w��g�a�
2��ÇvY♀����]�����8	�����Q�P؎�f'��W��#��8[��@��[�:(�P����cXHG�MDr���S�f�ǋ���0��ƑMBqr��*��"j��dz� ;ݺK��4!7��5��U8F3Q	�G%T"�w�R�|},a�����OC��}�ŷd�jrf��x�{���a=�FIQ���jSQJ��VW��.G��.�x� d���L�z7HI�牡7$��*Hg	��v�<Vz8�VҒ�K�qℯ�s,"=O��'aQ������v��@о���7� <�5Y֭�<(���e7�I�%س��)���]���UR3Y��(�pz�w�F�C��ڃ~���&-���[��X^�
r^BZ�'�}e'��O�^y�"5�%�}n�p�	���leʌ$e��<͙�����S:��2|=>@�������>m%;A������k'��n��w�>U ������,=��B��4�o�k��X����<�:*O���"@E�)|�E2O�R<��|ҳ$���_n#���6I�!�2k�mٳ)��gfB�@�%$�$Q�^��1�όՀ���'$�w������a��f�	�-�r����/~b����H�fOn\;�z-�j���xW݄g����Us?v����W3�O����qN�k[9?P�dB4���8�"7TV�����NM���-VZ�>�]�� ��1���UD�o$4 Ѣ؋�^9�j<>�����#�k��,��	s�#�1gP�Ƙ��i뼼���<�S�a����tV�%����l�n-h�$�Ֆ;�m<PK\J硸:P��V�ķXz��E�;a�)��	]�6I��j�[���!�gB	����Z����Ũc9Hsy�e��/�iD�y�HZTn��ݘ�rGy;v:Ӂ��-��^��O�5wH����Q�zNS��������OcK.��r�3O��Q�q�j6E���D i}�Zv?�=�Vte�[�ç�e�Կj�p}�i��<�b{e"�}�%aлz�ۭ�&��3$�|a"�$[��	G^Q�E�1�Ti2)Y094�
���]2$�[��?�#��-/�#%�<������>T��%��3[��Jr�2s�?Q� ��'���R�E���b	 ��طk�q�wߕtY��69{%t���a����`"��*�5.�[�ٜ��&��i�8��ɀ/�P[�������d���f�d�.5[����p����_�xY��)庠�@����OE��R*�"���\��#rZIq2O���f*����H5�:6n8����Y��r72V��ק{$=$Q~ѹ	��3�t����Э��6�����f��@<�Qt��;H;�U�n�}�W�۟��*1�_��5�Ex{p�ߨ��W�g�C� ���7KAy�z��6�(�Y�8o���� ��5��G��0�����t�7/I�!�M��>�T��K�d��G\�E/�R��*�=��9$�������lcl���M��X��N�b�SMթo�/���,7@��FBh�� ���0��Q �u���|l�{B�L���nF�KF�k�vLt�J���%S�;C���Ԯ���B4!p����ًvT�e��B�57C��#��G�$}{�xh4g{�ª7S��y��eq���e��Ai���uE�`S�W5mp��3��D��E)51�*�U��l��K��։���tȝ}ey���
��)�#Gƀ(`:7��T�6�:`<fgB�I�_뽯���}Lw��*li�%�g,��i�W���u>ntه�Ne���=��Ѳ����Q����$��)x�M�Xl�O�>	e�'�"��TrZ��k�h�UB�՜��j�v���iٶ�cD)i������|��Xm�}C)�b*y�T� %g�`���v���o V��v�os����~Y�qwأ�H�a2�S"n���4e�*.5H��wD�f�Vs���Ӝ�6OYn)��vK���e��k����l=.�[@~n�y�S���-U"��_��jh�Ey�g�S_��6���	�Ҭ��pf���GxV��3����� yķST/B<�oY�������Q,9� ̲�V	k��5�2��#�-U&U��ƽ��0��v��O5b�l��L1Q-�w ��Y��4���A�O��В憀�8z��S<�̋����q���~�%�Ɉ�Ȉ}�n�R��6|ଡ଼}ir��eik����ެ���I��1���Srr>�1C��@+?�3bJ��L(@�1R�z��J���q��rb/�y�����Z�Xy/x��Z���<R��?+�1b/j~��Ԗi��Zl6+2�Ē"�p��/����ǴOȻ7���.2iu���	u?7�
� *c��oRd�����v�K�1<���/�	y�Ҙ������m��f�����PG������m�<��֩W�3��ۼۧE�%���1��7Uf<m�z�u�wFR�A�T�Q�??��������!J�[�`]���p�c�pB��)�h���+��%��[jJڎ��"�D=9�%u���#�dNmǛ���"�!�uX��2߽H���s�j��h��ٕ�p5��6�`]�x��3vhZ1��5_�ѐ�5��O>��(a����Wˣ�X�-e;L�,>��S��| ZDz�4�m���&/���G'���~Q.����YǊ��#;E�p�$>�j�:G� ��.�'��_�ȈS߳ަ��0� GM�r�;RT�g����g��#�C64P��a4&k���l+��B���b�]5��0�d�f (�t�U���'̖�7%`�|���ݸ�y����R�{��ޜ�-�|�unY��o�!׭m��?G�"b��KO�ڔ�]j�����Y�m�����d��h���8����)X�{i�-w��j8��{ޘ��Ҩ]@�3����h�+���k�"�ư4n�Ѿl	.��h����f�%4&Z�U�K��i���HW������/�\�·D���2�?�lb�A�w��p?�dZ�/:����ۉ��~�<��$�S��ɔJ�d?��5����29K©�E���w��.gz:n�Q�E��d�&r��8n�%q�%jK��LA̪��Z��T��~-g�c`:3h�*d���E:kzNx���K2(
Ğ��q���]��(����֫����=���g��<g�ɒ��}C�qU�je�#K��&����.�u=��$��N�9wvJ6��ƚs� ��z#���mHr�����M��	T*$�����YK�e4�J���S����#����3��Ա�'v����^��Y(0t�C�<O=4�vE̿E���G�4�woi��K$f��9cI?�����D�p?����R�Q�1�AD�@���+��y)R"`��#%�|�k%o�tKC<�a�27�I{'�%�Z�ZL�R����XGl��Q���B�d��[�}:�j��W(�u ɓ��[׏HFG`�@��O����㼻����^<��@!w��W~0y�~������M5�8|�)'kt!lT{�Iǌ����?{��m���\�\����[�\��ښ�E��K�8�9� C��g2h�b�J�"ü�R�X��]�/V1���u�AH`��̧G���6��]ّ�[�2,I�L��ِS�b#m�����LuG@c�AsYb��#_�N���=�����E���k�=�<gTG�����P'��<����f��G����y�+�|�wp9P�i�����7hbv�86�!!��a#E?�x� �M ��z'�7�~�3g)�"����U����f�⇍�3�D�����\�EP9a��"�c�e��j��6�I+�vđxU��D�O� �y��7�dLx�u���'D3x]���yP��Y �E�@n�Y�G'lA��r���7�D�X8�|��S�G�K��u�~����~�WWr��*j��a��#��nb���4�K���aAν�'8+�8N�f"F��T�N	��_�,]=���+��]6�đ���y��(
��ɦ�o!�J��\n	=��M<XD �mu�q^J���(.1�m#�[�EV�+�Տc�i0/����'J"�+F17�&��ѻu͜�&�2n��_�v��z�^ņ'�L�<H	��7v+_5��»�c|�w�V�ؠ�t�y����]�}U��$B���V�U���jd���@�-�B��V�p?O�A�>�9j�몗0!��4�S����D��3�ݎ|Tũ
�\S(9�L�q�g�9���a��Ŀ�%�g�^��	=�8��@����flى��]��\�C�`���-pTc*�7 s |�&������.ڎ�4We��/�Ĳ��Ah�~(To���4��.d��D�|�����$Uv�2y�2ц(&N�������ͬZz"(�#�����l^ޫ4��s��m�Z2���͛ʃ�)�M�}�Y���?��VR�lp����B�/|�U[h�z�?e�M+��%G��ƶdV���C�^7���B��@Qj-�dWi�5����l& �PWwT�XK�j��~k��u��Z☇:�N59xf���d��L�\�����/@
�n<齎zˡ@�SG߁���l�k��S{�R�
�SÜ��Q=U�V?0�'��G0��UF�+�W��Ẋ*�wwGy�}�%m�+a��r>̚�z�=�3�%�Z��v���Y��p߭l	=��	<]җ��.EL#��br+j�s-D
��`9p�z���ڑ#�g<�r���7�y&��r�v
�`P��C�:�������l�������-<��=�U�ORפo�y=B����R�;BDx�I�Ff�*U�`�;>V��,q�.C�փ}��i�Ǆf�"6�뗷}��G?��>�s�M|�1��]	�Y�ǪP1G'[�Ӈe0 !nគ슣h(�.���0Yf�Y�d۳G|)�\�Ͻ���s�~�޸ܼ11��竈47	3OG�2�	׌����t���>|��/��i�7M�?��\�:�M�	>TH)�����������3.�!6M�Nͪ���pW�N�C��(H����'�n�V��3y:�Z��M�V��h�qT�4�`�U�'��b!-u,������Af���옌�J� �k���e4$�7o�%Ύ�ANaR��r�v�{#т��H5�P�'k�Km=��div��'0P�PF��םw�h,� C��ۑ|���'�0^I�"�Q>S.*��K��1
c��I�K�%L	l�q�Klc�<�X�D��lZ$а �DTg���K#"���Q"m©[Ծ�,B�5�bv(��~��G������M�2���A�#V *O%�A��u!���0�2	��-�nB�5�L���_��)�o}ꉇ�X?se���M!��ejOƸ����Eb�� ��84>��.1^2v��mnV� ��3��$��TJ8#�%�?��̩ťٵ4e���D�l+��ejB��hL���^|O��i�b� Q�ǧ���UY��+��9�4�+J��Ʉ|���
���55҄[*5�K�'�u�̣��J��̋ې��s��p}�?��׌lȈm'^![u� ���3���	�"|Y���E͌�gLH�+���k�{����\��{C���Ps (���x�^ʉ6K��ؑ�^�;~1�܉���v�P���qPnC�C���v����
���蠸Տyk��rPU�� �XX����;�%ܳ�f�r���^�^vFQ�u�O�����H5��{�*Ҵ��^��Q0˓+Q[���sZ����6=�F{U���f��`e��^�ڻ��qE��W���׾v:�6��R@��:3��FE�D�k����&��ņ��I��:c|�n@�R5���X}�rex+1hz���/�)�.�3� ��j��vR�jZ0|����n�mf*�{T��p��{Yv|���;��ֆ�+�L|�j�*�(6���uj\݀�,��i�����RyKI������9��b�vR�r�]�B��Rr{D��e<8�����h�� ��I:ί�h\��o��Ӷ���/^+d����XE�:��݉��(�vG�jؑ�5��
&��Qwf_����J�������`E{���^��?����v��-0y���Q�[�ͳ(ú�j��'�@�sKE( MS,G�bУH�^����B�����A]6"��v��TegF��?զ�shsYv�/4⶧ ���i����<{5����p}F�������9X�Ě�]��f$6�	-�ڟO,����/:,�D��50����}�/�(��h��Mew�'rzu���~6%~�+��7�L"�����BX�~SV��Y7�"�M�t�9����F ƶc��ڿ�o�rVf%i�m�M�����
TK�9�B}W:O�=5�DR��	�Ɇ6�ĩ���q�$�����6�B*�a����8�2�_g�Q�'ɤ!o(�FfI?�߮�����&��8?Ϝ��Sܡh�R-w�2N���+������C@Zųc�>6�bA�rk��x���)���
��A��$����۝��e�k}����"�,�_�0�b�4@��(G�⯲��e�;dO9�.�@��ޖц�����-I���+�y�D"h�>� ��e�8 �m����� �w�ؐ9�׎j�F�=5�Y �!ae��@Z�h��BPh�jGswy�N��y�bk�oV#dp��7L�WY��*��z[��<� ~�+8�y����^�l`-�ʙC��%��dށ�Mp�#�E����s�n�qK�̼e�Sy$xѳB��U�����j�AP�q!�s&��n�O�E*W�:ޏD�Xh��t*�e�^�M��c㤻.��t.N
�̩����U����[Ծ�<�ǯ�rÔ41o�2�ev�
9���&�Fm�s�lƈ���h02�G��'N��@�(o(h�����$l�\7�v�7-U��q;ɠ`��� ���Ik�nM��/>_���������7�~��4�`*�/�,�w�ofH�.�{j#y2ɕ�2^��?�C�d?"�x���u5A�(+��Fm0mp�M�'W�>�{��X=j���ބq�o�-�����|h*�	��c�e���y�x'+�������V�"l����<���5Ge^F!��d���C�$sA��l�d�2ņ�s�� U���7ɍ��Qy��;SNC���΁�`zq�y��j�R�ru�<`1��?����b���gؽ��'����}�T�v�q�o�X][7����������iØ�/ZZ���Et�V,�S��%���2��D�/t���
���^�p���H�D��ml�oRp�ޯ��Va���49kQ�DQ���?]Q�yv���'���|%����44Iu��d��8��d�~B��D���@})�_S4"R`
OL���(�);��j�QQ~���K@Ų�I�n�VvK,��,�P8^%�|�dH��
kéƥ%�W|�_&f�f��wx��X���c����G�|l��"�	��oE�:���V�.�2��جsI��>g��G��H����xn(��i�a��OT�tA��,�f�D�f^�N���d�
�!����S�JY�)�9K.\1�)v�	H��O8#�,_h���'���)�n�i_=�#��ije�q��a���9����J�OY�����-�v���<K��4K*�k�a|�������5�=§.������rE[!P�Znb���[�w޲�ܿ�`fyH��˖5��	�~��3hޗ&�g�А���߶ЖG�Ԯ����>����Z��K��F��)#�v�quy��k�qh`m�?�_����4A[�U����-e�~�7�eӰ���/m��:�����u[o�tJ7IK܇��B�w�����\���e]�Wath�BA�wUm�����sd ��q�薞(���s
��	��r�M%�F��Ͷ�o�����]�V�eM����Cd��9��z
�*rW���Vr�4��b����y�{����퉥�*���A=�#t0�����7!2������Ef50���f�W�/��d/��I�U�x]!qZ�%��O�ĩ�]g�:��>�d^w�PŽ�~�o��\l���ю�"�_���E�\}�[N'[<���|��^��<S��E����Μ��=yh>��s7�=`a����1�L��:	��ۛ7~	8g&����%)���uu�d�˝�w�f�-�^˔8ϓ��K�+�x
��L��G��(r�D�؏��T�!E>?%[<F�$��ѓ�����<+|�������W�c�0�3�牼�i��b�2,k(��(���S�C��{.6��J�/W~�g�����!6r�K��1�z�{l�ľ�S:+@��V�XV&�f��g��W��+�J���G�Y��T���^m\B�&�mM�>2�ԃo}�0Rj�歔���>��E��:m*Z��-ܵ*�%?���%M�3��fo�f%F`rm>��� țd��X����p�.�oF往 ��y���}2�[�Y.� ,�l�j��_B�[��5���I�X'kO+�C0��K�C����sf:A�'�6���$ȿۚA8+�D�,1�G9!�%=7̹ %e����7Tk BqM�ý�t�	2@�\4+{��9��/�P�Wc�G��T�	r005hnH�d�	��P�R3��>��BcO@Ȕ)+,w��=�L���6�P����/�������=AJ�~M.�a��!�����o$�a�&��N�kQ�]������E�w��r�}��k�}
����qA�a�x������s���N˥B�{�4���)-N$��=}�n�Y#�)e�����l�h��;���"M�Z A��_���}�1����WC���h�'�/[�[�B,xU�hOp��^� 8�h#I�8g�+���ɺ\��D^��aPbuJ �imuq�&�����U����w���kЪ��6��G: h�tC�����t�dG"	�cD�9�P�l��[ �� ?�	Y~�]�
���|��~籤N,��?ҍ�{���Ð����͚������R�\��>�c$�*!��V��k���W�p:?a^(G���?zтHh�D�k3�'3��"���Q���+��_����N!%�V��q���#|�A�ʫ���UFy&�<�d�l@�%k-y����8��>�B����ҕ��	pe �>���2jt�M�D�#)�u�Ǹ��
e��j��KX	��@�%E�k'��j���E7".`���N�F	�o�_ĭV���O��xn�t;&����Њ�<�nM��{l вN6���/���	p��P�����7y�H��З�۳fn��޼֎�E;�|=u����+i�����zv��%��_������a�
�O��~.�����È�\��eg����b�'0N��ˣ�L�&)��4239�̙�89�������B^f�8�ӗ������W�5r� `j-B>u�s��7�U�ʳ$�.��s"PD,�?�[)�RW�S����dkT47��C֏x���W�)X.��-��p�jMt��2��5g|ft�+X}���b��4�<
�f6)��?l��U��+��2�&�W�Д�$Uv3�Ed���8��}$�-�PB[��;�Y� �Ivκ�`Pj�HLY�jO-�!�1��� p|�=P���q -H@~��k� ��-3���-�F
7�~���ngBc��.��B����#����\f�03{�L"'+����#���*T+��E`�o+67��*�^���`�Ԗ��"� sA ��+J�*t�番��S�;W�_�G�5�@.�휫G��fz� �(1��1����L�������� ��{�I�LW��*�(H�N �|�z���h]�zO�[[
�AA��^�qQ(�K�9=������/���bd������4lYaĽo�'$���<=b��@.��ڻ��ߔ��D Y9�z@tG��7�@y��p �)/���2�v��p�ִ�|�Ӗ�+0���R��s����6� ���[=O�瑱X��C6CR���j*Še`��g)�_��_p��2�Ra,i���!g�
����[��%D����F��������WF��0���}]���?��q��,Wz���6Ÿ���]׽2ƶ��L�m�Ӄ�i���Ǩ]���2ޅq�rr��"E��3�:m�~Vr֜��'��������l.[��A�<0���2�'F��	��&�f�f��k�������vӜ��,Y���&I����ܐW>憒I<BO�G[�O������`"�9�k����b� �V�Ő ���jӔ��<zT��k� *h�����|��ǊD>�����ЪO��L�U�ڪ�#צ�1�7�����O��2��ЌE�v<�H�F�tMf)Fͺ�r�?)��Ixm�^c���3�(r��	8������B ���r�&-���H-�)2��9^�'ڵ�u ��H��mS�rf"�S�.�"��B�'*�Pw�&�^@N��7l9������R���X���c�~"�_�>�~h9�dnHg�斂��,r9�O�'yB9��8�$$mX�%P7 �rh3 F1�^;+�|���v]��
�zaT�w\F���\�6��Rn2dn)�>6�R߸*�hK{zC��<��&?��J�2�s�1%���b����#C�΁P�Mԭ���/���i��O����a?���*x![�fw��!�Ժ�¹F�&h����ŰD0�L8�*�f�1J�5�*�h�'��)v��tQ�֒��Y?���LC���|����-{O�����)��F�ݵ����(Ow�m#΂��gŻ[R�4�M�ZC��������lڛ��@����~�Ǧ�lUebU����J�ge������JbПN[(/Ǘ�I�ez�?9"!0.O[AqSɀq�z�)Yl)C��Ϡ�M%v�^�Ƒ)�=����;o��˲&TU]��垏H7�oQ��>C�ֲ�I�ΌN�.&��1Z�!��{��r�zrX��v�O��������FM��#8I�c�"z5�)�O��&�-Ѭ9[`�L_bh���{"�;��ho���L[�A�"��\J`�(jf�E�T1 �E���d�0����yu�ņ�<8���P@�en&���ۧ��_���o+��*w��q87~o��kQ��$¡�2��yjT�q���1��X˚���Ѯv֌禆�3y����a���tA!�}����\
�z���|>��n�u%|��
eS���=$�Z�%��6��*�|q�Z��&��B����ֿ��u���T��]��
_1�V#��p_1��H� jD�㌠�.9|\*�����a��"�<�S��f� ��l	z��`�ݗE6��K�����v8}c
�&0�/�!���1���e?�rd�~*�)�� ���,�U��S3�S�"���P���*=��)�q<r�앬���?�_)�sI����� �s*�wM�.����3�k���@q'],!}%l4�A��/�����������fZ)��j��nb����L)�hr�{�+�Cj'���,��Ny�u�A��n�pk�b�/.�e��P�ᘒ����_�`���j N��ބ�JA�W[��~���C��#��7���X���hal�?b�QU�6��{�\�7=hT�����\�:l�)������(�2ި#/���O�*8���ڷ%P��k<��I�do�w�:w��~�:���a�L�Y��Ʀ��>"�r>j�	H��
�_/��3����E��b�K������5[
P���B0��ň�/��\6�]�bl�T�A��k�w齾����u_�ȶ���y��;��t/��h�1�����E�L ���Y����Cd�Rb0u$�?�1H�mxV�7z�E�z�;�m��[������T/���H�!�:��%�=+� ��P��Q��,c�̛���A�RB�ց��*`s��YӧB$L$���+t���{_���?��p����>��f�&s�Ƭ���y|�~���La����ɥ�wB�E%vX�O���{8�$��FyVj��Q �f�0�ҁ�I
�w/�6%���:#�S=���1�o����vٻm�u�O(�c��aV�2�a`���H� ǫZ��W( 
��f̴f 3�+Q�{���v��	k�jշoR��X�����%u�9�(6���2�w똡<�[�z�OIn�q3��2�k�Ѱ��逌�� !QG�H+�٭�e�خ��Nd)�/��Xk�	�Z�(��o�hI%%����lV��_��t��;ȸ��T{�Pu�����*aP����^k;����� o�s 8�3�3�U']����A�v����2�k����P�ԟ���� Tx���m"�h]v�nj�)�× 
�0�ݟ����zn|v��\ߗ��{u��Y�@����R{�H�(�N�SHM���y���˅�1�-g?�*��S�?�T�-<	�������H�=Y��7��tB˳_=?��֋����S��%��紻��v'�5����S4����h ��
J�I��i�$���\Y�T�]ZtC��N���v�`=���8�ݑ]b!w,�u�$�>�
䙅�� ��i~�42�jpR.�-#�� �u�*�7�
���)���S?�M#P�Ho0��Y����.G�N�6)�(�j���F��_s]5(��r�)T�O���W*i���C⧽�Ko{�9M����M�B@nT�Z��|wöԢ~��eިM�@k�*9�"	g�m�x�����<gDy������������� �B�+L��4P�	������e� J�@�8��b�$�Ē��d�C�r��W�@�����y?��(��@���y�F��%!��0���b#��	Fc�P�T��p&R�Ҟ�|+��*�{uV�6t���m���D�W��A9��Ɵ_c���Hp�2��X����5q������,�S洊��Π�\0ݐ.9Z�4��M� 6�H�۞STc�3t�z`<�r�i�L>�����I��Jh��.os;��~��O�>�NK[��}^X�/[��]̃:����t��C�Қ��L�P�b]����ZU,�%����*�1�7to�X��g����ϐz���b�����U������W�����DW�;�|�0�S�<��S��ݛ[\�**�y�[;?�I����ˎ��ۆZGy�FZV���:v��O�^�����D DUzŹZ��N���e���ENCn��e0B�h+܍�%�e )���]�`Ϥr�۔�ؐ-�dE<c��`��r��f|:���e�s=���dn���]k8��i�\�z��N�\��@�|'�P���Ea�a�b9d2>�R��M�	��h	7�tc�4Ԯ:�1�����q�e�~X��fu6�U�C�}�M�����3�i�\���������3
k�`J��P�ȫ"N�/��!V
����,P@1��=j��:�����-��S*-�b���Z p����>�<��t��S��r�?&��'�J����N���û�_`Ɩ�i܆;;���,$9<�oY�d�KKI=��NZ��#�D�_�V��v��wW8,��_�|�;I�+���2�%�t#*C��Vk�B�Q��mÿ��-@~>��v�oK��>����N���2�blV�ޝ� ���W���&9�(�?�)po���~��9%w��GNN
�Bk����΂�?��Ū�*�|u��9�z��戆���^�:v��Ɗ��P�5L�R69$��3B��67���Q����ףh�|��2�nD3^N���x�D�X�p�iB�߶��a�r����ɺ�$��wcI')~��=���R��{u�
Q7ٴ'h�H��ӓ��j��f@��%4[�d�9�ô��{`��Y�������"�~�Y�L�4�	���A
���y�Bg{mű&�ڲ��?.��E�h�$�w���˺Jb�� �`�=�.k�hN�S7�3�$rC��ʣW��_Ȣ�xO�IӶ�l��}��}̀��G5톥^�e��=�T������mHk��23�
i����L�67�u;<O
�Ķ�>���H��VJJ�S�7���H���|#��k#��B��7Զgy��\���^(�p�X�
Sܯq�Ǯ�R����2+�\蘿���)Wc:=
eO����>�,�L
;������w�����$��3�Cd�n�ŋs�E|S���� 8�������hvKĀMUKŎb�F���n^ʻ�#^�H����ްҭ��yZ 6,#\J�i�=6Ӳ��ζ7{`y��pB{ϙ��f�8z)�e����ȷp W��};a���Af�81��I���Yc,k��	�������%���Q�1+����V�?2�P����H�So0-�B}���0��6~��2���
�A{���&Hm9|J�Z��ET��QD�5���g���;7[��{�u��kZ~�Q��z7W��3�ߪ�V����Ul*gr�=��t�ܷX�3p�W�֦b��[�����o���XB����72�R~���l4,-a��(��z�v�c�k"_W1�l��|�D���� s�9�|�*�������F�s��_Q���:F�mpk]�"�y�
��!��^����/`aP�k�q�F 9)P���\���� n;[�ш�� ���䯆5�ޡU��S���I���|�
Uc��-e��[Ǿ7V���F��曕�_���f��;9��8���e9�g;c2�M�h��RČ�v#!�eL���-��.~�m�mb�W�U��.�L�4��!$�x�&�#�6���Q(��K��`���˨7����	z�hmӶ���.yo��Y�c����t�0
��Bm�dso��t��#����D�K�\l����G%g�|��Y��!*��Q�6�\�T�f� o���{!��d$������Q8:۰��4y�%G�!�_w� ���#"����Iػ�c���O��q��R�C���Ĕ��}E���=���&�&RЋ��(����xJ�R=��38��_�h��7�D�c=`���?����-�q�D���_�TX�}�:R����쀟JC����!��R�����i-1���ۨՁZq[p��))<�;[���\���IUV:~�N%�1d�;�oې��~�;��P_�����V�%k��(�5D��Z��޿g+K�d�����,�f 9	���R�xL��u���s^�D�]lԢU1>��-X	s�ݚ�u�+z�����;�n�Q����w�"bJ��)kC�\�D	ԇ���y�1ٴb����V�!�3���+�`ꝇ�� ��~;*�$�9-�#4,k�<�6�V�UQTc����ttx�����e� ͼ�hԡ�	WP93C�1��uS�Ld��+Q��T]h��QF���w�!�+��E|��GY,�^8(Z�E�0y�
cJ�;lmWYhs�!�*��#!N�s���D ��X~�V�����TΗj;��ձ0��^j���w:�ǡ��W�	7�>T`�4���>��$�2hۃɇ��s\�/
u`&���������Ʊԏ��*c�Y�K1#����;mN��G5���H�qYb`s�1gkw_r�T>�1�"*.?w�"�|$7vL\<4U��@�����I�;R?6@Jg��g5r&��'��u�#�����N�	Xc5�(~�Q�;�����8�C�ʏ�kN�`��}�<n��_���x%E&�]�j�+��d�q5� ��� P3�� ��eϓ^ti�#���OT3���c�5e��f�gܿA���-��&��������'*kCiV�Z�2	�5�~��R}k���}m�%ek(���������In�p]@�N>�s��|��1d�BŽ�lBw#���;�νV�u�V�3)"��N�'�!t�_L#�Q[}l��6����l��D��贈`	�Qy��5�Z��-z�ȕ�Z�_v�����HzCG��G`Z�B�����3���fo����� /��
8�N�i�m��V�?�,��V+���W#~��P��?Y��R��o�Ð%dQ���y�2f�m���W~v��	�`��M9��:� �޷��x∫@�M8IЦ��q �I�e�^ћ�K�Ƹ}�4I����v(<�\��\[�^���
\�Ԁg�3P���٠p/D�C����u�]G��Pb��g��a�f��;��s1�L�-�}�|���Ԩ�<ʆ����j!��Z��b�+�n1�>|��ǁ��D���;_�b�l';y`�B]a��߉)�����ezN�l}T4q�s�|�GVǧ��VC�%W-Щ��3������r����� /�PrH%��d�̛�̠������+�	�'����ю��L���-/���
����2Ł��B�����A�D�L6n�����Y��!��`:���Ԕ��[fG1e��,�|�N;�h.�:����)�77tl���Xw5m_H~�E=ؕ�3�$��:@/({M��l�/�*gZ�W#�(�7/�Q�27 G�"hz�
&���I���f���΄~���fh��K
и�xԅλ[h�ABc���d�����U˺������`���!����רY��,[�|Ã��8��3����ʿP���y�C���4�����G<<��G���Y�c������jyֆ�,��8c�J�e�eY��ٰ��yR��R�P�h�&��!ńu��Ey�~�6�R��7k��q\Q_i��5�4�f�Zc�|Y���;��H���d��iL�+D!����v���jت�(x�����v!(��nbE��{I0-lt�Xi��+v��X>��DE��y�o�}Y_�C�Ⰴᇨ�@i5I���`�c_mga�r��ⷩ^�\U���0w�d=󀄭�0��V<��(�~4���U��X��Y�=���=I��'mU�xtՉ�;%��\[R��ZK�[25ӥ��@��VQ�B���܀��?w�U����m����jB t�@�=��I�o�"Iw46e�8�m�9��P�(f9`M�"�L����c�mޖ�㭡^.�翬��sy���eqU�Z�M�ӹ�ƽ�D�Z�t���\�'fy"x�e�w����j�u���*B���$5Q�:8����ڪ�H=��)�
���x��Ј`��Ql�*���F]2��lbbf�����R�%�ߌ45�X:��m(ru��5�ͻ�,F�^�fM�ۊb��.�咲��]����+��$)O$��H�2���$�VT�zi�����|.�R��;���[�mD��U�]��ݡ�x;zւ"��b»j@�#�T�,�ؕ�B��wMi&�����-�nǟ��*:��O�1D��N��Z�f��*6�۲�`���$���ˤq������!�|�d��H��tj�(�\� \M��^и�,L��Dذ|4�[|�n���x�Q:&!^>) z�8M'0']S=�.X�Ī�	��H��O�S+����m�/����50qT�%v"����W�&��_ݒwT�Sv�ے���/�6�.���q�_��� Fׄ����08#7�m��I�] �z_	�A+�9f�&k�����nVg*��EU��+�N���Z2�����h�����t�Ivu\$w����k��N`�1�{�������7{/D���GG����_&Y��������n8[���(��=ƊIt�=B����S�\�rVRAw����JttD���H��?c��=�2$%��~hF^XoAݦ�
�� �v*��y���:%�X�u\���P��'i<�-v��.�p��|�|�T���Y�� ���c�uS=x��JDN�ϲi��E�]C� �n��`f|_������$����s����Y�� ��޴��,G��}�HZ�1�wU�56wpH!�'�9���z�ͯ9�g聨d�(�y�-z�ʏ�٘_����&�����&	��Yv�F�%���Y�W��僤>m�t�Gz�*�M�ǎ�Y՝8 _��Ѓ�Fѕ+w��H%_�
���ڎ�H�_����/@������dV�2��5%Aq01�������2�y�bW
�^P*�h̺�O�9N�xg�~*$\[�Pb|�z�pP�/��xД�ڴ�2�����V��X��B�s�[޾����_��\%�S�bFՋ��|�]�G���b�|�&M��s����1؏	.�g���J���� �h�{�K2���4޲N�S5P�B�������KEÔKQ���R��@�R1��T)=��h'��su��0KS���?�B��]!o81�=���j���UI��l�׼Фk(_ʔ�+�Be���-��l��s�|��!���c���TKQ�A%7����y�P5�#����ua0~��`�L�i6��?�f֨�.(.i�<��NHS�wd&酽��B�öz��rY��V2�N�z��� �1(Qq�����U+6ނ��߳b"cҠ�>����?����'`��qd}q�}��@e���`s���T��ce*�m5�G����;����i�!�S�Z|�����h�`���@����r'O�9-�v�
���M�s�Q���e[iH�-�X��:6;�SŨ/Ie���A]#��\�{uT������*��ք7(��Ǆ���%#@�~���-�E� �����ʥn�-�����{��;�w��q{�
�"2�
y����mj�ܓEϯ��=ǉ/}���{�q�ų(ˣ.1m��GMP���)`9	_N�k>bUU
�I�N�6Kz??�Z#C[�p:�49�µMpm����( 9�{0 x'{ ����N�+�Q5~De� �U��;0��',g�`c;{��K�K�l_����N�ӕ�4�&R�Gj���g˷j,7G���sHǢ����ƶ�x#y�5��fT��F,i��zf	H�0ѹ��:{V�T�E |�5��C�];�]����EPr#8'����>c���-uɪ��?&dH���m��d(a�G_���r�G/d��f�[��.��U!�.����5:���m�j�A�8͠QuU��7�&^堓�C?NvP�0o��s%Ȯno��h*t]V=�\��M�g��&�'����-w�ײ�[�.R	�`�{x%b8�cb�+�7�T7츐�@𤿘�@K����p[}~�i��*���;H�S�/nʫ���>���W�_䓐kπRt2�f����jv�|Ml|��/O�D]��e�	�5������(Ͻ�0|̪�������SbgsEČt���#����	�9fg�����0x���I�>wX�ob�Hܧ���fR�q��h�e~�K^Md2�9K��r[^�I%7�R��b��ÿ)���0�}�U�Mݵ
-�V�ev�>!�~k�����p�q[Nb�P
ݢi�")��o�A~/�L��^V��>w��Ġ&嫈y�>�c3�vq�Je�m�m�C��[pL�F�&s�q�JR��)gWm�~ ��gZ#���{��5u��M��0� 7��Bq'҃��;� `>Ͻ�⼝�c]$�
%*}-̄"�����eȸ�;ݷ�͘�>���Rei��ޭ���|��\��'s2���`�UZd���qb��H�5�wX���*K :%���Y���F��xff��>�E�iOH�g�Tc/)n��+��nAG,��hpRAi��שa>��q?-XfkO�p�<UHٞ�6��g���dQ�<�r((��k����D�:xg�:��Q��)���-�ՋAa��~�w#�\f��F���x�!�m�$��'�N
�XVP��=y!GޘC��g��X�Te��2v=Z��������l�������p����ұ��wy�P���|�%��j��{��J(K�$EAQS#��W|N�ʺ�C~�]��V\J���v+^�����]�ꕖ���V��3����+�/����zo���TB���0%�$ϿK	S&0m�����m�}?f.�'o#�^�g͓�^�j8���ڎ�3Lz�mn�FV�"�]��Mrh�0����#E�c�;V`f��y���*ि�s	އ����3\Y�
���jB\��E/�bRLq 0��J��b�rj�H	۞�t<��uEc�J��R�,��.3�`B�	�k��1������Sፐq\�:3�=��m���^`#�����u�B�Dy^���1a��"�Y�&����~���g��@xE0��YCช�4�`A�Cwa;O��	�6&����S�q?O�y��2n��4���iV��p�N�gMu���T��A�h鰬X���%I K��'}�T��ئH�ͧa��-�Fۉ7�����Z�U�D���:�,[f���|7�S^����(8���^0���.ڿ�b���&,kg�J��}�:^�G�'~~~nA@��LD���q��j�؉��R��y���A��4��4��/���43ƳpTXv����?�+%�@�,^ꮧ�����e�Rj�2���jO����kd��}D�c����o�"�M���R��"XSԓT��u��'�L�����#B�QB,"��� #{B���28�Gc�0�ގ��K�W�9�\������`�	��zA s�|����2��bI)��۩�u.�i
|Z)���S��[� �|����{l�������c��,p
j2�]u�b�����%���� ݠW��\D&�gT7�2R���jyv"�F��yv帄��l��rd�kFF5�4��8�&+ʩ}1E�nq���z? �'�=��zS��PD��5m=�4`�0�5�4��&���Ozg3������H@<�·�H
w+K3 ���8G�F��4`/OU{a�5�7PN{���TI�9��r/�g3!IC��r�ʿ�_���p��K�����O`&�]lc�a�q�Ak�T�s�*Fkj��?� �ȱ%��%˥o$��T>dͳ�Hi����mO(cO��n� ���U@�gK��Ie}PN7/ mp�z�e�ΦQ�%mJ���g���v�vÛ{*Y0
��+��3zq�\�d�$�I@�'N�VoT�G-���{�p#_��x��(�«`zEBT�GO�H;��8@��e���(\�+�,�71�9�Ynh�]���G�k4ΥţTsJ�~~e����uh��In���Ԝ"~S�ȅhsK��^ ����:u�RM�w���x~�3s WiC���/Y�=���
@S�Isk��}�$�䭽�%9\�P�x˷"�|�����2fX�p�6���d�m��+�-��zS���6茠�%�i�L����U�|�h_zI֫#�������mF(5M8g�^����Q�����2�r��1������;�\�f-^4C�Y�����lI6�c۠0�@i���/��t�x��k���n�H�,U4��a&	A�~8���Pz���K���0���<�*A�;�O�~ͮo!�P�#�r�x���K�&%C1�2@lg�[P�'S*/Q�¬B���(�Iy�GE����Ac��|̗w13���C�`.���3�B0�V-=��S1�X��/���(@��$x�T�1����%�VN-���I?fnc�wle|{�2��C=j�E��H86�GO�C�B��q��P�7�K�W��cP�n�dͽ�jz��'..gAN�L�R����
b�����a�ſ��rh/��NL���<�ݮg�.$� a��J���2A�ؾ�@v�Qݎ'�жfd���iHdĥ����������(�Ӄ1�7���,i���ڼ"r�<os}�=X.�+k�Ƚ�Q6D�1�!����,��u)�1��0I�MV�'솼�$����
ގ�D�V�{�ھ�>x�\[;�^|��xԑ��6@O��k��aף1��Õ�*4�|ꎗf�|d��I�n�X>:ֿ�ToLr���Ku��AK8�0�H���8m�<���M,�ǎ�qbN�m(UQ��گ�dp.f�3���O'C*~� B�5,��"X\��Jo�.��[<)��e����I�`%V�)'a]Ւzo*Ɔ�P�I0>�Zu<Q�� y�'�Se��lii�����	�~dyz�ߊU����>{����Jڻ�a愼�7\����W��6����gT�ƞ)'{�PR���&��T����ǟzQ�7g�?�����L7����'�Ɩ�S��,����;)�4��=�Y~H�g��<��Ĕ'1��w� O��Nnݫ�=��Kav+���_,��ꡣ�4��)��*��Կ�6�uO�l����k0��f�lN�}�^�=����M��QSɉ31ø1�Y�1(;s�{�U�7~Jv��EM�U����aK	g�A��ut�-8$ӧntK^��6��S��,g�⒁l�G��~N.�B���`������ȅ�^pߩ�^-R_�{=�i�Z�>t�P��'a�>k�b�	��B�/�����y�	�D^����)�+,۵MǼ�ۏ�)�����\S�^�qve6�{
�R����-ü���qkTd�f��ǽ��:j� �%��	����w�$i�0�p8�~���)����\�m.�ڒ6��:.���Z�\��V�W���+ZLj�;h����'9�׼1���e�S��B�a4�_��_��1@d�6��x���PJ����%W5�{�Nd���6g�Sd����0k˝#�$o��#d��Xd��R�,��9�8j�sꎹP���w��l=a�2A(l��V5À��a��@�o�i�^2�>�(�'OgK��yd�'듀b�jX*�&xs�V�3l1�a	q`e�|;�h��+ȇKw�ϛVBB]�H�*�%=\h�'|XXH�7��U�C�a�=���A�wcHaj(�;UǱ�o�^��lB��O $�qM.���sTg�M�PW-g�{H#(��c��@�
�WG��hX9��O�5�R,(��OG�nؼ�>��:��Է-��G^��P�(����.c��{8|���Შ��G�ib��Ō-3�W�N$�3���|`�ׂ�*#$Uc�E.�%lلO���J�R#�XuV�{Xݡ!�������@B��a�8T�04�娖��}���^�n h�q'��J��n�(K9�q6�7�����px�:�WF���/���5�y�/�yT�=�f�4���ս�U��xl������N� X�.�p�ɕ�#'"����Jʇ��oՇ_�5�E�'�4_g�>^%�!���mG��+�H�q��R���-�`����a�v��>x*��ŭd	^����QV3v��d�g(�9$������{0��cӫ����Y]Nt5���
�Sl�������k���>��	�3~��i�����M�H/�h�.�!z_9� ��ǐ�����i���w�/q�\R�b�y5�\�B�J�g���äv^N��";<]�B�0hz��n�=˺sB늺�'�h�7��U����=,?'��,gv�c�T��$m�hBT�@��_ �r�8��� ��Ïdݧ�J��1�A1�;,��3���8�z��_=5�����g�~�#��E�UMC�dK�7���0xg���$�_sb��#2��$�g��u@��%e"N��I<C�7|ja=
�X��������ż�ߖt〇��_��Z�F�C����γ�J���T�#-�K
�O�;z��j��������L�!�f�e4��i�H��*[҈6��@.O<~�3>�χ�*��~]��c�<,���q�20�����|��rՍ�l�������K�Z�8�;&�̫�Úi �UǦ�gK1HאTC/-�4~�d?��~v�'����qa� ��������1FL9m�6/|�e/��YB���[��%��`��U�m�?�ޣ�M1��� ��h�+�@${�ҝ�Yl�1g��!�����R����;�rp~$��_�϶dF���_
'pe!M��Hq�T��	�n  �aj��s����P�FN΂I��0����YSD���o�(Ƀ:� ���7�Z1�H]0i��'9��x"n�6k( �5\\�Y�k��3��F�.����ǿu���i�/n�
�[�^��Ƥt63���f�a��o��K�"��x������+'P�������Jg)u%��i����:��M��t�	R#�^Y�{�n=�U��\��=�?��mƣ���G����ϭ����q�;(�����`|cl����N�\;��sq,��z1{,���m��{�/b�jHHjM�QF�'&=}Xg���k�A�D<�ɘ��Է[_r�/5wU�$N��h�b⽋/�Ȫh��5�]N�ԍ �XG7�"�N�E	ŀ�����xO��	�<S�'ñ�y?��'t���O�n��Է��s�N��o)g
��}u���8�J��%��*![P������pmb0�_m����JB��T-eҨ,���v�8N�H�|�?�htF��r��:l���Ƹ\����9�>��N��o��c�g+��U��®{`����-����:!\:��%��%��g�!G$��i�>������PRy��Ҝ����V�A}!��U^m���ޘ�LKלN�8���\y	�t8�Mǵ��͜�n�T���c�F%���I�g�P�� 4}Jb���'�,|��;�X�[�TtJAZࣀrj��n�װe|<��5��(�X�J��� ������[�sPq�2
қ�F7`��n~�AQb�v�b��:ՃE-��9C_}Q�F8�u�%p?v�yB,'�%��=��0{+�ZԔ�����Wg(���|��8��Cә\O��8���2�k�!H�8���v���
B���Y������fܓ�?��Ќ�Ԥc\�M _|l����Vi���/;ۍ��i�x�'����ǡ���	z,D�%-j|n﬌��g�9H)����m��.�XDF��_�q�� ګWO���ɒ��&/R%��fSV�n"������a�(�O��df��%p^���w�M�
��
��*����6�S~?�O�dϾh�E�z����\.�b헌\T�*�Č�f��	9�}H)��|@�E�#��#J<����3�ۼY'Iip���j�/��aH�L�b
�\s���D�w�	�3��G�}f�6\��4\��� �� �~3)J�I`h6���!�~o�Z!S�Ԙ��yu��㸆eQb*t�)H�o��)L�|����ܭJP���DM�Z�U�f,����f���[����n��%E��n�EYCp�w8����&H(���<�Ni�ti\���MB�w/o�֡!t�4�qx0��Am׫��Ѝϸ��ײ�E�=y�Y�b���p�hA���<� t��_V�2�>�:/���8F��Ȥa�Ui�}hq4"��˽�ע��4�Άg�2������-�K+ڍ�e5(�ӊ�@�Y{�1a�`6\ ��S�u7�g��W@P�d����M���J%��~Ȫj幅4�Kt]���Z+ʿ>�"�����\0��=�R��ڰ1�����杗�ݱ�=)�\��&}���mK�ߑ܈7E���n�� g�I�Շ���mjq�6����0�w�Pn(>[y�t*��n�5�MS��G��wN3�@��2�(�Nm�ĺe����@���R��5HI�.��}Hbu�������������P`� �U��Mq�� �bh�%���bN����`��I�+`�-s� έ�Nʕ$F(ؐ�������^��1�	�s0=b�� �N�5�o���7h���2"B�6X&�|��9�2C7���
�"����2��P�+L���r+��A�.a�.�٧�,���,�9~�>F8Ib�|���T55�3�\v�{�)5�i���:��:ĭ�A�?Qn��������ş�tOE���7���N�Lo�q:����3|�x p0�N����'�ز�"v��,��M(�˃Y��u���"63QC	�48\W-��j�=d8�O�Oj�T�q�-�g�I�:H���?m%HDW��7/ZP�oQ��s�w.Z:ն(@�b��3���M�`�h�s��%t��:�Z?�n�nL�]��Ƹ�'~���;,lEP\񦔟sc�o�Q�C���V}h4��la.
,����X�,b��Ջdki�6%^�����̎G]wV˿�17�"���l�t�I�K�m���qF���D�=������~:;�0L�.M�c��2h�Ec@}����wME���܆)}9o7)
B�� �OD��R�g89{ͩ��(߇��1�1̹���4-�8Wԩ����7�,���[�� ��aC�3~(Wr�@���X"�0;#n�� q4k����Pzh�_6�P�t�2�~PI��(إ�N���̬�M��{P�f>7q�@�e,��sH��
U ����S��'U��j�8;�}���ҽ�yȣ}��5�MH��n}�i=n�j\�@���j�6�u�
!�9������OBW���B�I��,xJ����l�8��W�R�_�@_���ձ�M�ҙ6D�l��&B�_֘�Ӱ���o"�w6���kE)��p�Ik̜K}H��'o�Ų�w�d��C[n'/
L��!%-O}8����bL�n����N�y�/��y��� PW���rn�E�IbX�{o����x��=��1�	l��K�U�	lt�շ��9c��\��dk?z�� W��4db/f���kL'��xG�O�]}�/���N� XSe�;T㟾N}��<<z�(_���L{4�c.��4]��*p;�Fdk*�Z�%�Օ��Oγ������ѐ�oX��.��Ӟ�M��fHi�ܔF2�+)�ѵW^*b�;/��P ���Jjg��#�H��Z+����-Kx����Q�T�^z97�z�mG��fϧj�%`Q6��u{��ܿB�M���bx'�^Y4h�@����~sFȣ��E"��*Ы�ucv��,�vW����U�#�Ug�
N�vr�"����z�%%�U�Ľv���:lA�90��dR�7��)W��¦;s����+���7�Q��9ͲR��c�*żV�`�1�cM)T�u���~�Du�W8S��n������z$I�,K��O����W=�4���dE3/���`��	�����Q8�ذp�����v�	ʆ;�`F�.?ˉ���x#+�Q)�\(����ܮ4�l}�7?N��(��� cC���g��T$G���\�R�˞ w[4v	7�5U͎h4���F�sᯅ�m`Ҕ�k�E?�:[��c� �pC�v��~f���jy��f`}�<-ɣp�u�-��j�V���Ч#lE�����s�ê,�������,^&����%�� A��&���uՑ��o!�ۚ���o>$K�L��fX�k��|B��x����B��45�C��t���i��J
�i]p}�2d�F����w�[�ۄ�������5l�;�Ǝ*@=�]0����=�!��t�cq���Aغ���տ@S�H���j`�֊���X���P�ʿ�382�=�V���$�i��b��k�Y�G�EvXރ�u�L�`�� DC����w�$y{����e�H�8�>���E�H�O�)�,M���>3g��܀�#�aèY�a����g��'k�E[���8�sY��W��	��n���9̗|�88�a����[�y��o�b|��l�$L9o�:Ľs��6n�7 ��d&к�6���DNL�~�gԲ-}W����)������ږ�sz'G��,���L������h}N������Ț�)E�
�P�}��F�D���Þq��(���� �����u�b� ���?4��=����S�7y�n{�zeU ]���J�wc�{��G�y����
{�@P`C��jU~�n҄L��h�oD�˩ė�������z�i�J�p�ĭN"�O�<�!����镐�X�e�u�M�[�t�����fT�@��X�á�!�\A����Hl.�*�Qr[��@R�%�"�#dqFڇ�%ڢ��3�HƖ�F�~/>��&SŎ�fÐqO7�0P]�U|��#y�����KG�_�|�!�BM0�w�w��i�3&�p�<U�pড&�����	�e����z@�-fˍ��T�ap�;�<�-fIIY�t?������X�����Ҧ��=!"���E��
���?au��ϴ��w}ll�K��[���-�j[ |vS/d�u���0#�(����45��n���]0[����*�8�d�//�8����Ḁ�.�H�,����J�;aqh��!d�g~Pr�2�#d��x5������ȱ�k��G�Gx�}��3gBN��.	�AG���IW*�S�����@���r$���?�f`�X����gX̛��ˏ��= ���~�[(zh)�<�I�<�G�zeXҬ�>UG�
��v�)���8�e�nj����I�B��|�#�z��i�Á"x��u���R�����<��%���yJp#��Q�F�*��.�4��Fk��?�BT@��F��+N�2O5t�B��A>��%�b�Br�-� ^gz�� �L
m��>����4�M޻�_���bh�� �:)9����.)����jt&�QVI��,{��G�J���
�E����}_����(nx6�WEQ� ������@q�^N@x����$��s�9	~ݴ���ӷp����ӚY,FL{vQ���*ڢ�}<�[��]��6����lP���]L�X!ǚr�.�67ĝ�O<����>��&�Ne|uG��|�6��IB��ec���N��	kt#�!�|}i5��>�
����>��h�m�L���U�j5�J�����D���0�>����f~��6O�vm3(Q��>�����z�X;�d}��
�:xm"��=�f���V�ǜ�%�v�R�&�g5��qen�_�,!0/�Ob����HmgR���+��;�$��k�H�dV6Q��ᔕ�Aҫۖ�K��6�����u�qꋟ�z�	��Q#:[��i ��uӧm9h�w.<c���^d�I���s���y^IԅZ��ES�
�d�˘W�m��t.��3Ȑ� 7l�� ���W���
����#��i��E󪪓x&�W��޿wH��s��O���p���2�h��:8H���ğ�
�S�;8�?��՚tBAN8�}��!�qe A���h�ݿ5��Ÿ���XS�.�	�gZ`�ոF�x8U�����S_�
.�/���W��:@�
yVZ�=^bͤ�)	W�1O�\$?�l����T�����>���9��]_�$ V��(�d���=d���M�I�+U���d������-��`.1^Ƶ��G�L|�>�������>GV]���x�G��"j����7nv*R&�b��=�D):�>�oRޥ������Sɍmn4��3��m�x���.�oZ���!��9���k,R�.;�q��ɹw��CAA/�A,a*��B�H,�},:\^��?_�{���1�o	E-�Ϛ��Y2�
�;h�~�p]st���+���M>7�b���sO^��$�b��n4/:�S��4�V~���\�*�~u�Pg��L��V��W{�L��~ �M��hҶ��4��Rrl���_�=R��j�k��>�C����L�BP�~��u|�" C�
���щ�?�08Z�D�+�p\DzR6NVt���
�4�Œ���G�̱S~��0B����z�'���;7a#��K�ￔȉ�j���9��%�7i�:JI���B$�ੑ/zѻ���_����>q � �\��~}��.���8���?��ib��<Y� ��U������嘘�9����&�]OC����f�a5����poP5ڪI)���D#%���y�G�ᆈ 	��n'���2;)��>-�����X>k*���j}��bW�=uP��q?��pV��}$m�Ǵ^)}�_�c��y�Ĉ?�ὡ��r�Ќ��>[1dq�&F]��*6BEhۉ\!��S��{�Ds���%���H����)F�ɜ������/�v�~�V,NrQ �Hg�u7��5(��Wр/�Ж��H��پ�<f��R��1g�<\�4f a�G��yd�oOGk��Mx�#��;>��6y�u���vks(�;�zY����i7޹��dnkOٖV
H*V�j��L����Q@����;iף\�$(�96�|�k(AY�+j��m&u����ZE%����k��!_��\K�٢O�N` ��@)���C��f��^%��E���X�{��\�v�"�?@ڇ���Lg��V�5c!��Ǫ\�_�,?^�Wx�(�*��a�w�ϒ�,�@�CT��`�PaĦ}�d���p9	 0�;��:�!9��,�G 3r�u�SQ�ɼ�I���� G^����AƇU�?$H��g9ƨ&�~̰}�)�BG���	�R=�D��.�:=�DK	��&���­��9U��\�p����֝d۠� �n�L�p~��Z��KA�m
E��k�q�* v�v7���xL��HD�v�:�FZ��3��܏������Z��Y�̰?yb7�J(vJ!�)�C��V�|�a�h��`&(7��l�h�Sf�O���9VQ��C�u�^D�
>"�cp��ZZ��?�L���v1�n���I�-��Ke]Voոw2x�_W��d �E��$����ۙ��$�J�4�ӡ
r4�"W�4�<�l8����2�s�#�t�Ͼ��3qZ���RӪ�Q��BFx��A��C%{�br#̝v��"�!ś~Ko��LA9�X�����j� >���*f�շ�[��O?�N�t5خ�߲��~�ۉ�t9[�G�1vU�nL�1�a$O���|�o��W	��s��J̙���1�㳸�rK�LpO��,pu��Ld�w�|f1k��+I��o6�{�n��X� ��
��f/6p}�ڔ��Q7��˷�ʻ1���&����y�+�L�ʄb��}HC3`ZM~��F7p���`(ߔP�Y��R|���#����`�ە:$��j:�� ���26_?ha�It��*����y)!}�jm����ê$�T�{�C�����י!6�rh�f�*���e��%���.v���lK��_A�<YVd!E&6O�9ʊs{��eN��"���K�����VB 8,�I��I}<J��r�'�5Z'�����/#���g^�ai+F�U�^.EǭJ��ɚ��Af2��d�V�:^���[BcV?�����ʕ�Of�V8Z�Q��S�+Z���9q�hN`gYi�ľ:�N��nD�{�	�@��p+�-��}:V��T���H�-uS�Ln�.������Y#z�/[?0�A"Նd��jA�T,��3�c^HQ>���Į�Q�����O�og�9p��3,m]�r�"+��eV#�?�=�4�����NP׍�?��mH�e�<e��l%�����߄� "�z.!n%���1����vm~B����Z����&��e�;Fg.pE����J>�o�T�Qc ���*=�\�SQ��������i)G���dm�оw֋-����柤��ۡT��Le�	|ЍuY.���{��7M�
����8BJ��s�k��f-G�e��)�j�boΓ�F|Q��{��Qm��je#���p�]����*k���H�v�`�9�(�9{0��A�����ܖ����c/4��N?׭ l���^ݡ&�N5`Q�Uaˮ�ּ��C~ �Y�JQѬ��vF/���ϔI�-	���͛���xq�u!+����9녕՗���C<��,T �#r'i�:����p���G�(��>�8~S68�_�@0g�������A��ޛ_��Hh��C�fvQ���ۃ0��;;�<&[�
 js�4���A�#�;).3�aY�K��w1�8�.ת�~��>�l������2�3}_/ԕ�� d�\���,y~�c�|j�7����9@�ʐ����7�%HQo�g2�8�el���Uy�M�%n;f|8~�PP�2���X���D��ր����7�g�|�h����+h<nj�\3�����q�XRT����L��||s{�P���z3��W����LȊ��&�Aq5��'��e�('�hX�dX�N����r�}j�[����F���2��;�Q s
$f�|���8�zj�ȵ��^%+�&�`�<��J����W*Q�99��!�9��悔�:��f.��{�5f3?84���F��t ?x�a�L�/��p��!�#�M[����(7��D�_KK�R�����]�&��YK-�f&`y���wt��!�}jm���?�7v��D�!��r�@� �bE�ǉƿp��bޓL�X��|�:ռ�S��. �_���V�E�.kF9�i[��N�-A[QlM_ ���*�jZ��")Lq����;g��Zq�v
���F��щ?�_�s�l����Tf��xKx���wt���=�S2�\o �O_.��;	��`F�b��:��'6�Eڲ8�f8X�?��s���G�Cɍ�*7�J�%4��cTމ���b���5���R����>���hu7�i�L�0n3��h���T�]�lm�T-��{3Etcd͙µ��d��=���*�N��Kl\C��E���9<Y�x`�9y$Ό�t��Z��N��Lh�{�����RA&G��ddD�p�lS���Mt�	,�������1�tX��x"5������cb>�=�FY���pZdΒ�*#o�MwY.,p��}#�wI�����T���3;1^x�a�f]A����މ-3��	�46yݛ�V���~V�?�Q7X�5F�6�=���V��k'�2���)'/�רo��)~���0���L�s#��c0��ԱӮ2켻_���ղ�4A�ݪ��iH�=\w�	����,L��ڷ���#Đ;���*3U�����1)g���m׎X�b9r��G	TGdFj���_�x����o�7��Im�@�HNp_����	%U����i��:(���s�������J�ܠ�a�Ps��~��v�T��՛�U/&R�/\�}��1�e��_�>v�%[?�r�e��D�uK2+D���H�
�� �����Fg5K�]�y�����4��(��ʿU�ua�yz8%p��+�M�2S7��d������1Pҷ,Ad�7a�Ϭ��[6gBMa������]�m���T>�<�c�s�F�n�h�$�Rf������|�VP@�ʠ�%U��g�\q(��Қ�"`������V �h����e�0�0P���J�:{K���B��.�N5���s����-��JP;�_�jɷ�eE���/�&�������	�2R�ʙRJ�'�]t]�
�GcyaN�����_Q�z�٨�8�e5�d���X*��w#�v�C$�z����|�Q�������Ge&����#��8�z��ȺW��^�(l�KW��p���]0����' l#��>�_3��١���F�H��w[e-:}��1��m�\����ҥ��Vj���+��l](�}5,���u%D��6d[5/�c�J��w\F!��K�' 2��
M�e�����G�A���i��I��~lL�G�h��s���P�S���Rmu�B�����|��Dw�Z��'v���r��ǝ3u;�R������㕁���Ag�ߧ���.6$;��' 9���ϯ����Gڢ'	�m�d��R֗�-�#$؎P��bi���@�>�Kzu���AS���B�iY�C����)P4�Z�o,&�d�Լբ���jv��V��w�*�f��n�x�!=��2`����(�B<]�w7��U��RwqF���[��
�=we�
�Ql����',%척�e"F�l�,�1�Y�[�n�tH�k��
J*�����m�fb���.
���+q"e���Ys�Vz2gO�s�F-�F�
8�B���!I��4�d��Y����6��Y�:��/��B[m�T+��%ȯ{X�R6"ے��Яz�a�e�(�#���&N-~�2q�t��椎���C�����FU' Q+�8Ԅ��o��eU����&�uӠ��-=?[�N��>�a�9�GLD ��$G�2V׾Ӟ&�,�g�A�)����+�lַ���d��0�74+��ެ+�,y�8/��Z����_��o:�-���mIPKz(Ǣ��� ���Rz�2��!.��9y��{�s���qsnW�H�����n�9�dޤ�v��|���)�TUk�y'��9b���lit��Һ:���e2��e�]����E�`�I�ܭoP�^�|�3��g�9Ȝ��G�%*W/|Ҟ�ǈxr R�Nm�M[4��H�v�H�E���x��Ao�^#��xa��r�j����T!w��Q%Qt�}L��g
f�@�MN�^F�	\�����j�����E��9�6��KG��T*�QA�]�tU�q?eoե�֑V�R��
��G�Cq�s�{�1��E���!%��j�&���*t.\6��%����FA��`�ln'-�s�b��{C��L�Ү�J6j/�/�Y�(Y�ҵJA�7�5�7ʺ��Ot�����,w�)��ݚh�V�[��}��7��O�Ʈ8��4'v��-X*��2qG�=��������J�z����{�-f��]��?��д0ϺW��� ����C��c�,�Y~�@�4�J�@�^pi�P����YɪCg;�L���R��9m=�%D�����7�O��~#-��
�׈=�Č>���)�Sn{���O��!��ߐc��nM�^	>��Eb/@B���&�ȚC�D՞�����'���Ws��+��%q���$,��d�o�s����,L��~uSJ�}���g �#r��`�޾@O,����g�n~!rmd���L�u����ACU	��rc�_9TxZQj	!��.S�;k�vǻ��7��g �s���K7�L���5�j|LMM�a��VIP��.�H3,��7��ѧ�!q��� �e��<ٽ���ZT�N����n���tE��u`P�*6(�
`�̲j���d���۽rD#�؏��,�:�J+"�g/�G�U|�|��$��s��73}#����׵�c�:�;�;c��>N%�D�m���]���s"��]}���t%ȳG=aee������|u`�,Jpz�w"$͜��.of�z��~{_�W``�Oռ��UK>mj��l*�
��?��K�+���S�6�38���x�RzX|Y�J��ޔXM��#�`J��z�o�8�n:���1�;j@�ïOx�a�C�iM�~��m�ԿL��`5�U�f-�ƙ����q3X��E�G_|cn�B���m���fX���
��Z�v��s?�<3��_���Ϧ�#��̣#���	^=���Ӑw� [�%԰}��ŽÂI��o�����W������]s�ܷ���[٭h{�jp<�X&y�~�ըdt�n>�9��s���~j;Co��0W�`�G'�{�� ��]��E%�_N�Z4s�Bl�s�˦�3|�u�rH��"$�� ����C��Ƃ��y+�+�g.Y*˔�Q_}}�\�le~��E��k��؁��g�Dʿd�֐��ə�t	��\�Ynp��C,>$���x)$BA�,R名I_!�󴡙�b���X�}�K�6�x���&����S�M�M��Ӷ��zd{�t�"�d�>���,�ɳ�k�m#!��й�d��;�?R�
�ҵ��e�c����Af1D֕_5\��>�CQ�1�����U6��}��Nb��KS��ګp-��&�<6���)|�TvCn3EH!�em�N^P��P&�����g�V�?�}�Kˇ�m���y�K/ w�RB&�l7���Am���e��:DA�efY��X�ƹ�}�YGuD�QC���A�/���V���a�d<�}ďT̸dEj �����^�R~�{OV�� 9�A Z�.�픝�Nϐ=�[;��kf��3D�TqK�a���B��BT
+�Od�,$�3���a���� �T>���3*�. ��W����g<��F�(���I�ؔj8���$�!R�@;(�~�̢Ma����kE/d2wd�i#�E�f9��٣��g���蠂6��8b�x��v�f���	�_-N�1Es����d�A9�@TҥѬ�]�X}�z��� ���z� ��;+ݯu��|ȄٱTkU {�rZ�q"�FM���j��;�NHN���n˹��m�z�"�N���R(:��~Q��ql�:H�n2)�Å��zUW8Wݨ�S�]٦�A�����|1M+��)ù&ChBܲ5�q@6SL|K���;�W�����XԞ�.h~��u�|M6-�[^P����c����@�p	6ʪ�U��%s,�m�C?���&:����3��r��ޮ�aK5L,�I��/�;�Z�i�I5R 4%�#��&�[KBA[�y��{a�i��fV�s ˲���V��xj�Wh�iܾU���f/�M���B'>/��H��+�>`Y�}
IZ��)�ȵ�p���f�N)g0J!mZ0����&l��:3�;sd�^�B ��3#@�����B�[)�=S�.�aU�>�g$�:x!��Y��W����ب��� ���\��fA�|H���nߛaA{�_&�1c,�{6:���nA©�Bcl��G�^U�/�D�ZQ(#-� �y5(9��4߇n�@n���Վ詎*Љe�$��Y*D�6�~�-nז7F�^/�l:�M���H_=�ņWtS>�k����{|�o)2���g��^0�����"�{,����K�L�'?{d�:8i7�;��/� ��-�A��j�F�f�?�5�ȯ(��qə;>z�Q�����7	�~�֌&���Z�ģZ�<�� ��I���B�_�逶@��RYg������d9���c�����.�c�V_�)����:���Ĵ�����1͠�ܺ0�d̴,Q��Ұ����]-r}���x3%�BG����q�o��5D�ฎ�.nc��0 ����:�#�c�p�s�c7:J������O,�� ��؈G�c�%�p75Duў�V�ǦMo�ݸ~�;����) �
��4v������*L)�a�'����c«��r��5!�<���C(�a���wIrD,��;��S�F����f��N�6� -Z��H�!����<�W$?�<�,��-*$���ٲ�O�*�+W��<�i�\���L��z %�~n+f� �������r��zF�з��G�0���������s(3����X�Bg�ȕ&�.��e(<�������I`&��v���S�x^�r��	�Fg)�p������w�oź\�ֽ�=�Hd"�$p�����_&8��ѓu(�($C�& �H�|� �*��{�˕F��CtBG�#��L�\ŁAD<����A�D�=�����Z�An�_T}�Q�u����Ulw�Jgn��u�)�߶g2e�w� ԄxZ��&�y�`o~K�[�ɦ����sV�r2��u|sI���y\ܚuMF_�[�uӤ("&G��������E��fzc�ܪ�}qA�s�Swb�(�O�0�'e�c|���hG���xv��w�s�_Z��'31�e�<�4*M~��u����YI���L���QxD��8�
3cu_�]vuH�S2���B���8FܶZk��a&i�����}��9�"J�w��=�t����CDO�.$8{	88տ����+����:���숲������ʶ��Q�D���ٜ(!q�CS�_�SEc-�^�\�˾>�dm�����OP��:��ZH�Pk`w����¯�>�+t�g�96m�OJ�������m\$n�k AP��z��a���l�;��/�����xo�2?�ذ��q��',�Ȯ��U&[(#�sB8�D0�V����eʧD鮟�m�JP�[A��̞5�PCf�a�B��O�M+�����W�/~-��&'���J��ǔ���Q����<��
~|��P��}Ց)؁
7���&�۬�>��ʱ"�29il,B=!�Z#�S[u@k0�|��z���U,:=N��]'�(D�{b��Q�����6~��g�ع��h��8�ߣ�%~ h�V���t�l��>O2�4ai� Ae6�Z%^�&!6���J�%B<��I���yu����2*���;�D��`ʊ��l=5�4�_f��wَ'�P$;F_q��n���.5F�{�	�}m5��x�uiƸ�ԤL,k �v1<B�r��.�Ҩ|k"P�!�o؟;[����J�`;��j�pe�`E�[:���gR�@![!]p�~�����j���9�A�ѲҔ&j5?1sM���G�P:����1.[-V�jyM8u�+ʖZep��ܲ`��+d�y�HÇ�ObY�/��9�p�J�-N��̎`��%�{���L��B�X�Ϡ��k	��b8��<��OZ�~���ZɅဃ0g�#���g�V�4�Os����p�𫺿pK���3%�IĆd�Ȼ�9}�<U uZ���R�W��HN�x���_
'�Q���.=f��qdAy�Z��I��r�U��G]q�yg�@���������}�@ПNWs��i�sE�'f+ꕏ�A���|l�ݽ���̕~2�Ġ&���=|<�.1�m�9+x1،�J��c$a|s9 `���8�t�w}�ʞp>�*]�f�������zT�R��ƃ������sc�|ډ����D��-��_��|�'e(���zu����]��/ؓ��ޤ�̢TXW8������?�вښ�(2�p)�8<�Lo�5��U)��0�Y��ϗ���vo/��#�F��g�R���ߧ�L�� !U�Q%,-����]�;s4	o����\g��Ev���x��:�E�X�Y�X�wP���z�H���C��ٳ�+>�#��)�7��=�K:"�FG>��5xd��e$!D�psI��X�i񄥡&�)���*��E7*�fB���`���Ǉ���o3,$���]�xpZ��������i���P�d��VW��윫~R�,���!��T~w��d �R�)i�.�Nh��ǟnM�eع��IH-����FW�;��۪ߤ�j�*љ�{%Z��N o�ˤ ��)�ۿ�w��y�a���ь/���R��b|z	�6։@m�VEv��ٷ��jk`z�t�.���l3`����R����l�k�l�vp�@�h�SHV�����E.9;��a��-c�'{�{�LS]Czû����#����T�L����(��F�&EHw������kP`p��b#� E�0l<P�����mhq�R�8&pqq��I��9- �J�%���	{�cKx���-hZ3��O�;?a�H�������G+�b2X;Ci��b'Y��@=�Yf�W��P���%��;Q�
���F�@D8T��~)�X, �wO��h7�hb��Ja�����}&(�8Z���x�=y�S��0��o�t���w'$��&5M��V�4_cA��6��
WތO� �ר�SO��1v�X�sׄ��E�������?Y���;V��^Z1;=^����`a���h���2�E!,o	��n�ǹߝ��o��	��#n���@L'ߌ�5N�z o�K��8zx�?��7�rT(�l��*�e#����Nl/�,����*u�@�r�d�� ��S����������-
�P#��u�Jy!{��X9�ێ���� �6��4��bR�'�њ2h��S�������k�^���˗׻�WUu���	�S�ё*�V8 p5���zz;�Pix]<G�YGgߌ���l-�}P;�NPD��d������p޿|�w{�:�.�f/T&�LZ3�	��5�n����i3�
�/Zs6�/�]=�g�BԪo��ڼ�ʮw�N��U���5u��u�Y"���W ��©qxJ��fZ>���N�期���+]Oq>�Y<w1��Ҹה��L|6�e����@I\�����6��Q��2H��F;B5t�P�X�g��7����r�
?�|Ron]�J�:���o�ݍ�)c~\�5�=(�X�c乔a���FǾ���yvN��g�ѷc��c�5z�켱{�w�W�ӘA5�A!�!"�ֹ�W𝡼dԶ\�R�W�>E�7q���a{�  z���3�ع�x{�-�ĩ	�.Y��]�:�9�k/���F6�m��+/���M�\�w��<o�@Q^du�������#V�>
��J���^9_1px���Le��&>��S�iYq=-e'�I�^��;�N"��į�i7��}�SP)�7DP�bwr~'B�J���@�)�h5��$���VA�࢞�l֒�5��e�t�-p��n�t���z`~ƳR֒9�tӃ ݪL�ɧ�@�6	�ݱP)�}~#����Z<+�	�m1ڹl�ˉ}K2V���f{�<^_'����� �&��abW��B�^�{g��t[����A�t�������m[�Goځ���S>P�`$ص��7`�vZ8���,�U��/�����#?irm��k��������m���}֌���_��f�\�\�u� �kAv�x�r^{<4�C���h�'�x��F�Q�20'1q�/y2�%��Q.���[U���{� G������@�_H�x/�&`v���4j�2�ĺ��
�����Fφ��ݳ�+�pz��^&���[P�ꞟ��F)�c�� �n�n���iG����'�B�r�Z��dv=&7����xz�*ǧ����xo�n���}08"����~����.)[��"�ۤ�� A��^/�\J x;-)2iaBNYE��8�U�<�g����t ����L;����52f`N���4��VwU�=�G��ؐe�G���O0�=z�ٜM)d�^U�'��<�k ����ȘPL�nTS�ɉ
j��t���%_3�G@�.�u�p���*Lx��9Qt8�#eu����u�T4�� aѾ����%�l�wJa��/,�S����_�n���#v/�H�I��}��R�q6�mQ2Z�<R_xې?U��q�9��yq`JR�dV�ҭ�(�z�RӁ(����CF���s��Vf\��+@�?�2�ȹIi�ŝ���	���������2�]<�[��u��	��F:d~�eo����{��νވ�9�6e�_�mFe�>�x����N{�)�+��R��K	��W�Aq�ڹ}�+��Nvs��h"��y��h��~o=��fa>�&�q��$&��Տ�r��v<���W�c��30~�Q��^mM�.B��,���E 8]:���ԉ�0����N���<_J�U��1|�R��O�;��M�?@g�a��#؊,���?M0Y�մ�,��ʂ��F�$n�e��w ���Skfx��>�
�|J�9�a��r�50چ��Z�V�YAl�e��}n����G��/|ͽT$Fk�J���߇tZ��Tx�.��w�_.��
2�9�B�=<=�/��}AB5��)C-7	�����P���m�����X�\"�
�-WB�z��1&^c`n�[�rLIIoŦ��1Ouy�4�bG�S��OLr��_P~'�Y�)W�d��u\,k}�V���q�
)�Fη�p���!���c��A�`�ѩ^��{ba�q�jt��ʀ%��J������-p��6�ގ+�2���$hކ����=ԙz稹;���%m)��3�ٮ�;��7�GyYQ�j3y��Xd&�D�,ߏǲ)�|xV�&I��R�m�M�mV�
����+�>W��_\$^Z��ʨ�"î�4I���2!v�NA#9�l�Et�e���_Ï��z���< P�;j���]��%_^t~�>5�-ClY���)��6��^�h�8��&�h��Cv�V��0�˛F���UB��HM��!t�?�&b�-i�4�;c*D��&��'<[��+���d @���f��D��|��2#Fߗ�����إH��Z������E]�
�����)3}p6��@�z3�Y�^�q]
x3.~Je�T�e��惬L_���ɤ�)N���[o��9u~��� �U�)�[�P��y�6/��"Zgd��f<�*A�>A&c'I�"��K��e��ia	�L�b�O����ǫ�|ez�)�}ic}�:ui����%�����媬̊�<ye�X .���ޅTc��˽����Jf�#m$����ɉw���JùV{<
�KT�"��8Ln�u��5�~���nmJ��Lu�(���� �]�5���@J~��S��c��-��hK@ru��� ��%$9Z|<І_��cC��(E@�[�Y^�& ������D�.��Oܛ6��I�l�s�x1)E�;WdtW�i�=ۙ4)�h���d^��#Qyk��Bk�#��:�m�!f1���à�)cl<*���:ē]�m]�Ag��[1'�z|��T������!���{��x� ��/��Z%��˹׷�S��8t��;���!52����[cTr�O�����f�����C�[n��?���%����)1�jm��ኰ�$zP���	}4�:���������en��֫��y��'�v(�@`�Gr4� C����M�9�k�]����4������L��z;���5|�6�<� 95��%���_���~l�d�A��l:ψ����ly�A�H�!nc��C�R6n3��͒'��}J�;��#�X_:^L�
�7y�47�s�$�G^rW6^�j��O�dux�&Y��&����,^��ʟm�~.�am�	��sH�au_0��wO�f�KqǼQ��V*�?{|��B|�<���oS?)��z�����h"�9J��1�o�Q��Ǌ�b�D�������1��EB��)�0�����@j�vŅ��<-ʴ	7F iVZ�P��eqZ$K�e��]�\���ǿ��5��y��,mMiul�u)�qR嵭��c& M�Ě@>����4�e輊���h߬J�h�I���W.<�J��<��=�dz��]�K��fR��d��%�<d�
lCJ����e�T`v?����`�T����_�/��܏��u�)z��h��We�����P�髅b�C��*"�A�<!��+"���9$�h�c��T�s��r�qS����>+�/�����K*��;�5�8Bⲵ�P�{�LQqԧ
�Q�g�b�;<휧�OkV��/�|a׻)w8����U��lI!�ʠ?��C�ó�$d6�G��D��i���,��J��R�$~��"�����ۋ@�%�� ���D ��ۡ���02Ryo����b;lKɒ�L��φ-�<`�� �c�ӷ���&���|�[CUH�e�(���,��;��l�yY[�8F1u�roJ��p�i�� 2)ܽ�q����a�ZXk&jMx�TQQ��[�1|Z�r��rH�9�`�uV�L_F���Sӱ���=ޫ��#@�߸���C"��-ke(���`�,�l��)��
>�u�/�`�~,���kgO��TƮ_�DQs�.lW��6���[H[xPq�:M�vPdB�qжI�|��$��|3�s]x{�s�ĭM�;
��ۈh�B}{l�������=8�=��`�]F��G�ëhb�C��!xk�I���
GёB�\�6��+���o�i��X���/�T�hjk�QB�;7���D$|؊3�kX�5��I��!���7� t�t?�y}S�;��|8�9�*�@	0�4�r�~�-� �nj�a!��9�5`5�姪�Y^��xN \1�81Yi�X�kJw��al�rl����4��0����R��T@C#��l��E�6��j{�8¼G�����O��F{��4뻕=4��.���A�!��C�fv�ȳ�_�o��> nb귿��Ћ_�8�G�!�(�
~/�a���y���Ű�~�:���0�kz��� u:vb�ǠC\ɉrw�q�)$���y�q�M#r���r�qf>�o�����- ��
�T����{�7��,~5�Hh��]��0��'VT5/ԗ>��7�-D�܊���&�1`T���>fE���3��%c=B�V&��.B�Bw��i���A	�#���ez���$���vi)��<0�l�ηU�N8������T�.��$������>�����p4Es8��Ϳ�Y�#�����s�N��~�-<�4�'\���OEX��'��w?�#�m�>��WI`�^1|z#�x06U�~�*fɁ���BOǽ+[雛|$���V�Dh��J�[��;��l%���@�?J��Ñ����A�4��wS��P��B~%<����h?���ENx��p���5Nf]��@��t2�N Q���������tCg�O41g>O�ܔbЌH��&�-��}')�9g�J�<���F����y�.����Hw�W_2~�>�+�K�j��V�̋���%�x�C�<���|x��?oZf�=�L6��v@�G�\�����t���r׫F1�r�2S�t��Us�3Ȫ�����Fۆx�_k��U�Vox�
�%9��N+6��~r�%�#��
�����V����"s��Xv��c�R\kжF�����ϟ!Zq�$� 	�����Y*YQ��c9Nu4龈��&va�w���f��d�P��K�ݠp�}'����|PB�!gh�<�vX�l���`� Bo�v/N��{ͷ�'j�Fq��&�B"�N6�N��Wjh���O-�"EIC�ż�}��nx ��J���7;9 ߶��E�3���N�������)��)��� �Q��}�.�:e�D�\q�����GX �O�÷��	�S����Z<�Ha�UꛫW��y�$���M-=�wy�3��0��y]�]�پ@ �n:}uRnҦh�J"�L������ʴ���l+Sz��:��=��D��Eq%�
�ݻ��Qe��cC:� fE�7�\(�Ϲq��Y�uK	U����ɚ�����u�<��	�������sЧ�һ�~{/ϣk�h�R��)b=�����(]�|��8(IbeqR���+Dd��R&�Y�P�9{���(y��a�^�o��&�^@P*MI 
/,ş����>��C��ܾ�A�c�b$��o7,:,�����Je棕	~�za'��'=F���z�C�t7�fӵ�?�=��<K��+*�;�RK�:�"�kھgK�U�T!���9M^����F�w�H\���,�-�-��}���
$��5VQ�p��ә�8���jb����x���B�jke��nΰ�%FE�t�)x�����}��
�xM�n1��H>�k&��M�g��}1Z�l��?f\$1�q������$��\u������
l"�:�g�������|�����ҲV0��@'��r����7�ۂR�s�T�E�l�
�i}?���̘S��a~��.�E�_�[������Ԁ*n3�SI���rIq^�,'?&pײL�ԙH=tFl\�+�m��u0��åy�?������l��x��d�Y�wH�� ���v�p�`3���iQ1�#��*Ac��f�%��~�UeE@D�'�.q |b0��#��+@�9@ ����G�l�*�
����E��p�e���V�����c�'p(�%e���C�8:+܀�H���/tћ�5aٙ��M��LY��q��B���e0�ތ��<H@�i��~tm���YX_^���2���}�h��| ���d�^����w^�����d���0�6Ե�iϼ@?6}�C�j5-�}
�Ī�WO�E��s�-�d�h��,�g��e\�R�B7!�eU�Np+V�l�Lj�d�^��!A�e���<m"X���G��uw����u�.�c{U��ȼj���ű�q H�U,6��a|���s�(:��5
��;�sܗ����Sځ��hF�����SG܈�Ͼ�߈O�u2Ѕ�ܘ�H�b;Z��S��Ы�g���E�j�J�2�l�/>��k�h������	;�����>w���ˍ���w<D.����nmʏG!�e���;1��Y�_�m�R$ ���vϪ?͸7&�c���;�o�f<�Tq�&4%Ũ������!!W�<�n򑎿�1�`*1�������(筫���Q 2)� �ק�lm���`p�����UC��7R�ɕ�*g+'���(ɰوF�n/4��);R�]:�.�U*S�X�=;��p�`�ƽ�iE@T�� 3M4{��*s�*��G�������]���pv�0���غ��*�NH7S:�񹮋�+�j2*�9}��gF����ݾ	�o�(z��7ӱ�7�f�y�&(&�~äZ���̍�A�~����R���9:�2������do
e �h����*PB��FF)Z�d�-3N�1˸�DۛdKC��B��Em��NZ��R�b�
CԒE���j��kMe�{I`��Z��D~�:Uļ\:'-��p��#�A>��:����>VCÚQ<!��UH%?�C�w'���
�������hx�����������c� oHҪ�Zy���J�/6�8���+��s�%��a�Kb!��1:[��\a'�t9:���aq����Ǜ����@�w���MTKB�9��|D��t���09�b�+��<w�8O��a|��p� ���9Ȃ	a��i�]�����n�K,�<`C!���g䗅�]t,��J8ժt��i���}�s64Sڱ�j(j?g���j��� ������i_V�]R���聅�+nJ��|�6�a0���,t%����j���]��V�0�2�
�*�ɧEL`5" 3�{\Z�J�T DFN��/+��*��F����\$�wĂ�a�F~'��ʴh �������2�CW>��D�<,|��
<�}V���J�'Qgʨ�s�7{�bd���>rܥ�XνF��AO^O����{�|ܲp�.sm�
��il��6�	Pi�d*�hl��oS3����A x<�GP�e�E՟]d���:��W�d�u��6u�]͓�IK�(BKGA�4����K��v��G�ܘ�&��F�E��սMJ/���Y.�j�l^�ʹ0�&U*�,j���O�ɳ�x�z���q.��8�Fj�s�uq+�h �S/�*\���<A�E&�ɤ�s��m��eH��2�kԒg��.����pњ��nmA�tg���]Tfe{�{1VM�<&�o����%K=fGڴ�1�]�ݐ��W�8���М�<z�rDK�A��Ey�*�Ӷ���&�U��_�G�J�����O��p�+������� t��,���@��^�$���R�P\w�&�CSco`��W-��M���!S<��z�e8U#�&��'�M�
��PJ�B~���63\�<��@���6�Y�M2'7d^Q�Jh�3'4�o�|(��\[�����Ϧ�I_���{�V]]�m#2�g)J�Iw��i(�\� 
>j�F��e��wr| �ElMe�+Ƅ��C-��b��l�u�Im>LV���Hڐ�L�{�,��
��9qK�(
��H�g��G01��<�NnG1X��:}	i���KB��9��{��%6�|[�-��ghto����[�1�V�Z�L�CK�T�)E �n���T3(iN����� D��E�X�y�_���N���w�B?M�\_0bP���}+8Ͼ��^ �SQ�v�@�W�W�U�#͇lb�T������O�`Y� �'�Pf�`�����E�����--���h@��0�����G�#f�_I�$�uN�)��!����kp�g3�Y)[�vRwPeA�����@�.�Q%طZ=���qx�+t� \�@�*�ݭR�R��j6�ӫ:)πӋ6X}(`�Ƀ�M�Ѯ�W\K��)��vz��O˱t�p"#T8�A}RxM�E�nFQPX��k�P@�d#i�$O���;�h]`��I���m�ø�3p��E��D%ڸ4$.1Z�z��ܺS��A�O�����q�f:�z1��~�������m������<g%�t�)�n}L:��IoT���A��s��w��ݒ� T"7q�G��M���B���w��u��U� I&帷/�ct�Q	/�,�e���r�Vt|3�VDG<P��Y-9
�A�L!<�=A{�Y_U���:� ����%ߒȻ�M� ���Ƿu�e�-��ǽ|�� Nb�h��Fա8fJ�:J"��&����3F�Dwj���҇��Vx+����~��K��l��!O�oqCkV�#-xҠ`a�[��^�{+b+�#k�y�,;�Ms�G�.k�.||�4�g����I^��/Bh4C��Q�x��w@^���'�wgQj�E�g�݆�R�d;ˠ"A0զݚS�xݿ����b���^n⡩��\^P@1$�����cQ�I3gteW�(x&�2���0��W�]˵g����Þ[���������l����R5���w�g<b��ne{PY$^�`E�HJ�+^� ��rjF3xУ�*e_?� ם~���uT�W��\��NE\gj@a1>팠���"������F�U>�� ��_۵L�	����6Ou�d㔦�x0<o0�*]��9)W��sAb�O��0*,�D ��_�Oc_��Z�N��ն-е��_��\�ȣ�Z~�g��>�4��?+l!8B���L���ʣ+R������Ii������5$�}���~s7 �v�MB�j�*C�5��f�?�u�>GL�SO����8��%q����6���J���j��o��㚲U��Ք�0�' P��D��N����ڳ^��i'x�e&������`A;�0qB�פ:��C�5�QW��y�����bC���Yۨ�2/�+���d�o�«� lC�K�����Kj��ŮN,)�Π���2���=G��E*��M�9��g�d7�&�T����᫟�=��J��V�&�`s����S�MR�5)�o&�n	���N�*�h ����I��h�A�p<�S��;��T�L� wƱ+8��lm�q{'b��~�*��=���3�A�M�p�?����3�b��WZ����Âu���Z��߄�(�����7
�T\���k��!��L�f�\�w_b]L��[�'-�T|�'ɼt�ڱ�Uay�|��.�B����B!�E�h�)0��p�d�X���F�%.��{9�/��/��{���z�q$��:��t����D����Z��	q06:����@�g&�N"X�b',
?�����.�c�?��F#t�r��h��i�t2����Eh�|`�����aJ/u@��E���f(CUDgb8.��~�I��(�E�=�W��ʍ�������D��W{�������@��E	�?Ur�e��>��X�l�n"�����&�B:�� ���o��\�<�f���i���$wӼ[�}��-Z�|�C�?�X"n�8C�ڽ��C�q��#9��YͶ�4�Hu\l�+���d(H��G.���ٚ�dR��kS�JG�5xbf��Tt>���R�1�F:���!0h8=�~`ϛe��x��9�-@�Cep��0��u藔{�*ҡ.�]�ߟ�o���A���hfڂ���3��Q9��Rh�Is>E�"���\�jeЏ�������g_��h���y�J-�B$�l�U �a
����~��"M��{���n�h��7��|N�n��ҽ�ϭI��;{��ӆ�.�����#�
#���t��-7��rH����\�|���� �V-'�I��� ���u%�\_`��ȼ��^o��%�͸|W4����D���m�P1�SJ�KIUb�*Cq\ԚE�2Q�'ne�n��|���ck��_CM՘+ʸ�w�tZ+5� ����;�3̠��F3�x*�		�~\m��M���[Gr�$�3�?�����Q���ǒ�%��>�c!4D=�"8K_���mu�MC)e�'G膵��7��\���}�I9 �iw.ɑw)S���������nذ��Q���Zܿ�*\�G�2kB��J�B��HD�qv"Vv�cm�z�h���|�3��t��=���5i!�%�5s�z�� �\��PK|���\��!�w~�2ܽ���_�J�>7R��{>$�^9H�F��-���h�R8C{(ʕ}����wHz)�Bj~������ux���/���O�<�� ��RjB�&K�l���W�7'Տ�ve�-3���I�BSGn�d��ٻFn6)�I��@��K\FB�gJh��m摒�#j�}�L�{����T��ո%�ֲl����m7+T}�?��3?��{�ep=�E1�@Go�-v�"UǄ����q �_�9���C&�\���TkW\����)ߘ��*�%<WC�f����qG
"\�Ȇ$ɒ��D�,XW���%?(~���ԵC5v2���Ql7�<��g<|o�-�i*p�8��[Ὣ۶��(E��=`�4��JbG8�!S����R����Iݺ5���\�/�حE�;+�n72B�f��2rq�g%xz�8f��t+�J� ������Ø�L/���.\�M�/�[q�G|! ޢ-���H�o����Z�y`W�Kӟ�D�m�< ^��Ĥ[����`�r�׫��պ�\��#��/u�Y}�9�?�1}Ȳ\Y#��;u���D;6Fi�6[=������Ů;�v$r��G���И]���[�ZK�"���N��~�i�]�*ߩw�l���u|�S�f�D��Xg7K�@(2��uГ@��L�tl~UmM6$����u�;M�wF�[��B~p���'�Hx�F�RGX`���%LxOW�:�;I�xӀ0��o3�����/d�?�?lYo�(7�q�}�L^7�W7q��C��Rk
�y��P]9x�)HG����U?�ɼW��̾�I���{�>o?��?"��퀌&<������EH4ZRzMARV�o�����b����|�l,{)P�˹81"���F���W�2�V.�y��nk�����n�90e�ܑ��`����q�e��b|�. 3�6#��.�3��J�6�e��7�E�yn���%�.�O�_�#9��\~/�������M��f%���M��pV��UM��-֓�9x�g���o6��S�ޯ��^_e>��\�'.�0	��'�j�)~T	������w��AF�9{�+��0�jga6L@|��KA�b�v� �����4�f�5��+%wu]����*h����h|^���D_Xba��b("�g[N�ǋ�L!k�O>i���&�BD߶�9��`�����y�F��z�N����,V0SO��RV�yL��-����Ͽ�m�p����k��k�V ^[�@��v�e�N��F:�}�R2E;q���sf��or��'�S�fo�oLv�%Yf<0O�yp��˒/�1�[�"��,��4\��IQkt�|���! �Z��e�a�����梕}?��2CX����g���kL�TK#��F\RF{�R1��m��pJ9C�j����T�]r����(�5S@E� 8�Qy|H�m����#���+���Q��s��6�����4��O:��J%����=����[3��O_!���:u�/�.�
x�R�%�I��1!Y�R�4�px݁�� Ⱦ�@@b�6�'�-s/28͢��A���?UN��V4b�{�^HA���x�TD�~�����`��%�Ǖ�m���t�n+ܶ����s�9$\@Qu�ĳ~�bKݍ�"D���oG�t�Zx3�TqrC������r㝴�6�yp�D`��mSW�:2`W�o�봳!#��0�ݯ垧�!��R���|<��g�.��;2~ǰ`�3�Ro�3�U�Z{�+�j]��X�{I"���v%�ţ4��Ɔ�^�P��X�������Q����R�N�k)$Ӄb>�W&q0I:����BB�3�|����Ҭ��T(�߽�M�W9ed`��^m���.��vf�����}��E�~�30W9Ķ�U3����rt�3.���&7�s3�)�E��]�M*ʬ0���)��(ɺX� C&�qB�w'G�ARc�:�O�c��xxx�u1�z{q]5�D,=�s��m"jG������|8�I���|t(��[7*��Z.A�(�e�>��o�G���b�= Cy��+SH���E��y�����C¿*6�:�4n�}���wC�[cc�9�u�Ks
�>U�&��.����'�(�b�h�F���[px��y?ZU�$@(��k�uD�^��.Uw^��=��y��=ĥ=n��������T�aIZ�n3�Q׻ �$ޘ�����u�VM��ꗷ.���tMF_��U!Y��+�֜�����ߒ�}I&��l�گp�������.u�0����'���`&"ŋr��bC �S�L*�l������DA��c�I�����8*?&�t���:R��]��T���b���_ڴ��E�.$�u(��X��gϷ�'3�祠⭋������m���Q�b����o�'��=2�'P�������\m��zr�â#U�|�VYTgMK�����8�]3���9|JmA���T�%���/~�iӱ៭玥R��>� +���օ��@3�(�y�8ͪ������lF0��:D��pI����i�cz�7 �s�ylS�'�(�V���=��X��%�*d;�J@���d��2�&�"�s!\A�q줺�9���;q|������||3HgM3��f^jX�~Ԑ�i�ۣ�9�jwM��9�?ª=��0/������[���qkDI�[2����~�WZ��X�lF�>��G?�K�X�F�k�����O�1P�Խ�"-�y�R:���9��l"�M92`�t�V�e4C����>�@Hcc��G2	R�w�g+�A#���'�$Xj͘1`��l\�U�}A�_^��BC�	Äox��Mp�V��o<Q���.�"z'��/(�$A�����i���sNk!ʁ�6��-��q]1H�k�i\�Y��5��F�m�{e�4�\��(6��F_�����E�r=�傇oJ����Y"jo+&��ަq
U�HG�]n2�\��h�?c~�%�����(3��F�?�d��u�q6���S��JM�5��o�&�T�}��=�UT�Q���$�;f�3{�j�i�yvJJ��t!��K�ˡ`�U(�@���#D�q��ޣd�ulv8��l����D�����������iWD��"�K����+=�?we���&����I�8[?��C����j�����c!"SM����߮F�d�{J����1��d��4���������G���޾�ѯ�����{�g�W�?��Q��u�����Ħ�{� ��<��[�R/�t��+��de�5^�CB�u�n�	6F��O?51���]xʂx_1ݹjxg�+�� �]E�B�P����+"�H]h�H�[;#��m�;&f|ϸ#)�XN*�(B����$
U90��,^� �x%��*�X���Cs1���6����2���ySn�I�����̷.N�%قy۠XI�d``�1�C�Ef�0�^�ݽ�N�o���t��4|0�T�e��	�{
���*�Cݢs�3�y�&Oe��L�K*�4��-c�)��u}��]�B�8Ͳ�6���6����p�v^�2\p�dK[<���9o����*��A#\�a䧸`���i��U.�0�������R��*���[)n�Z��7@�]$92j�ц|g6W��4:Y�_^3]��&!��E�5q��'����;,��I�����%{_�����9���,J�wTK��j�7�z#3�*3�R}��@�êuqF��Σg����3�r[At����n���l�Nx��Y��g��Q���	J��3���s��$�Z3L�x��,�H&�Bh'jRq� K��6T��݋yG 
�$=!�e��;�J��p���(㤿��#[�~]��ݖЌ��*D5s�<f!~3�+#���Y�Kb��N�B�]�X�q=l������ ����Or�~@{�lz�2�J�*L�bG��+gq��]џ��`��%���d�ܠ56���g��>;P�ʭ���4�����W:$�qN�	Y�Z|?h8z��D��^�IPy�A�O���դ��������r�5��d�B�5�amq. q3U�����k�^�U���m����hX��rQ]�1r�3I�����5G��&��/�剠�u�2��+�ɠܪj���T���e�hl�W�<����sH���4%�uV��Ys	8K4#4�PYh1�V�����8>��١�s]kN�Van�1%���f4�`>��C�;�b��͸�hz���5��탍=�`��Ry]0�p{��c��R��������]�ѯ�c�;NwkuI�L����@s���L��1�]9��T;��O�A�&&��-��0Ma+�����h&��L��R�H�%�J���(j�'6Z]��e����������r�ͽC[��:Z0�����(�f�h[���� ����r:[�
�x;�券��Y	=�=�s=S���y�-z���0��eY���dJM���C���:���q4�-`1Q�q)_��$TWLB�h�)_s�D���B<�L�$��>�vD��fWS�X�w�D#�!�X����7H{�����D�t|%�)��vK-��?a�n�%_@`vZ��w��^	�3|�}���Y�"1���Hh4m-��-��m0��e &��.-�Uȕ�-c�@:G7��B5ՇeL|�$��%6��hw@R7ŀ=s26�h��˥n�6W���e�&j�����t�_�pG�0qW�b�(�[��k��lnx(p�����4��u����S�~�0��U�齐�Q���|�z��n\�=�,p(/�D�t9�YH���F����#Ք�(�����B�6����;P�u��N��δ�dS0�A�zf#Rv	�Y-lY"��贍�$� <u��`b�Ve�-KFڙ0?�]���l�~A&��滥)��Sw#����g����qy�\Ae��,��9�)o�$@$��HS?g^��\�� �1?�����p��T͝t�@��*��f��V���(��C�n��ݟ���_�flR���T���t6�/�� ˥���6G b͍��:�6�`L�U�c}�\�>���+��a
�.z��R��9�����P��!�v�&�O�;p�(�U�I��Ԉ.��⁥��/���q7��G��}���U	BIeC	�@'m��3Y;���JUU �39�$��:P@�~�ʞ(O|��Yh�ĝBEi�Ά��м����0'�E��������kS�Z!Z=�c@����u5���'����_�~��_�*�QpI����#{R�M�E[)w���7��R�mlB��ߘi-��ފO��(nv���B.N�)>KM���_�h�< f`�����_��"�p�����=�ZJ�n��~m��Q&rŰ����+VwaH�+��\P������oA_Qs������`�Υ�����.��լ�q����C���;�@�8��t��re�{�&p�� +M��7��W������*�����)���<���T�w�pu��-�>�f&Q�eo�8XY�r"���+(?ؖ�w�tX9[�Gc$:t;:���b��|蒏��M�>��x/�f
X�z�?�k3|�����N�R���cn�����AQDwN��+�|
�p�7!ʎ�����Z �,
�A�4���u��:�����[�4��	z("�	���O:��I_}��2���>��G�C�X�||�[ ?�������,������E%O�v��N�c��p�l��5����,Γ2d9�M��QYh�����[w�Յ��������#�,�iup���~af(��5�?���h���ګ,��_|�ox�`�c\S�����MHY�������Z[^)"8�
��4�:O�_1�=����2_9�]'}�����E�7R���U���G���%^b��'@d���mq�I�#�s�6@������<cKG �����ߓ���sm�-�d�^r4�7���s%Z� ������+5p�-ICPl�߿G��܏�O�+ȝ7����p��!�e�ن�[�L�
�)1M��P��� &�lq���Qv�h��?����j��Xвp(�$z��6|�&�.t��O4~��e��������k� "�c���$#e�o�KUX&%(��MN�4�q�f�gHkF��q���I�.��^Z|Z���P���<YRC��xk3��	,����u4O�ք�3��^���YЄ�H��^Lj�g��M�V�^�[��f]��Qr��!�� ��P29��mn�%^5�Y˸ZB�[?�H���8���A������.�Wl���xzi�]��A���81�C����G��x��e'6�rE�z���Tᄐ�{����]�'�j�_�(�7�8
�Ϋ$�����Z��0����O�Ay��k�e��3g�L��^��B�ݺ�|��W���o���կ���N�<���2{��j����l F�S��Ͻ����L
��H���X�3�����n��|���T�6�g
��Z�\�6(z%��*G���w�?�������L^�+�?H�rIr�_���E��'���Y�{�ȇ(cL ��N���~S�pn
O�4�(���]�b��$V���$��1�+�-S�U�bo�5����s]
�+��(Gr�.k����2P��qA��E��H@||��#�S�'r�����Q����i��AF�I#�Q�=k����J��4
����Е3�~��Q?l�Y ���y�I)|��5O�8d�\zSA]ڥ�"������M5/�%�0#j��S<�@� 1{�ާ�-�E͝�e���Ko�^�Q��3x�|X�z��Si?�K2�N�����~Q>�#	Yl}Ȫ~{9��bT횅�����Jg"���e�kID�K�YTdʗq��LK
�:�hDf�����i"��oI�a�[����,��?�����dL(�+���(S�5�j��=܏��(����|2��j�.��XiA�[�d��+<���6�>�a��䚚�V�@_���B��0Sq��p��JF��#MR�Y+�\nI#�ɫ_Ҧ���H5�R~�� U���EMz��3C���̴Q�We�k��v&�K��>�,�!�M��������B����J4|P�b�	�D���r�R��mmi��	�z�<Mr���o���7龱Tc+�#�`A� �������
hFF�V>5���D�!�+~�t���!��>AH:XP�����g�d8T�;�RX6_�W�:\�J�_�ݟ��N�~J/;��_A����-��!QR֘;ʞ ' UҰ�f7�6��Ɓ�4`�]W����.�]`�4X���Ǳ��(�����4�:�m�J�7 7D�~�#����!r�0��E(��
m8�ռNk��Cl�6=&$ ��|�u-SWu9�8��w�7SMcQ�W�;��H�] }�r��/�p�c�An./��E~����Z»R�_�r�:`�"�W�?�RU(�h�@��/�u̫��|���ΣL���{|H���C�O�LB��i��WE�`[������ n%U��#��%J��x�K��ϊ\b/gޫe���FY���ˍB����0O�C��ycd_��mst��d������^�$>���9W/��CqA����o'��5\�s�}`l)�##4�����&���w��(�x������m�b>y!���?��"ɸ�<��[��kǇ:��̕p�׫������`�@�?��ɖ3e����	U��̳L떷�PqaEulAӋ��,q����5#�X�7�k��T����d8���o��W��XB;�%���9H�l쭱o�?�ܥ�������zp%���G����o?��Vm���>�YI��r���>7�(r/�U���_C�T��]�ޗ$r�%��'l�k~��m�)�,xJ@���ݬ���"]��]sC�y��aN�С��`| y�*����`��s�,�"0����}l���e@aҰA}� M��=h�������ʀ��.8��� 7�3Ccx
�!ь/w��&&B��S���/Fo}S�"YG��k�D�a�����$R�p�e_< }�]C����%�2��b���c�C�*���Q�)ujRI9X������&�7�˷�^���lk����Ɛ�"c�6�@�r�#�� ��#��q������sa��H����2RѺ�Z6<l��[C�L��
�ʺ��L�e3˨N	\i��V�& �$��X�1Ϻ`F����O6�my�������I��j0���|<��&;k�`|
���P�*w�Je@��&��b�J�/r���q%����I~�?�o�E6���C�*1�Qy��)c�V}R�-7�j��g�Q��eU`���2h\g��:��O0n���婶SQ(A���YƟD��F��WUg�2��M�v>�� 3��9E*02c�1��f%@���'D�)э
؈Xv���x.�|Ѥp󟤥���Mߞ�CC���ә�Ɋ3Tɀ����Kpv�Y8�ʙ��|�e�+:�T�kbyR̓C ��0i����]́ǆ/ �o���wypRM���ݑƒ������뼷���bǸq�����H�ɚu'P���c�y�Wu�l��9i���(=�(=0�<���JT5�����c: �"[���]���tUXYǗ3�N^-�$��8B����<&\�b�>�'i�;���$�*�;���h ��������İA���1|f�)dⅫ�0����]4���˘��=� T���O��E�L�C��7핎�1]T�xс<�_d���@e���9���isV��m{윝��u;@��9��2��h�>ʶ���D��7��w���X�C ��0yb�*\�J���%P��h4�S޽��f��j�A��R�c�8����ꃇ���ff�y�*�tȜtQG�|L��n�w�b�?V���}�o��i�5���>aT�,�1)Z�PeIt��p���燠�D��M�c� �V�氻3 �q�>�H���?y����7�]� q��{ �yܱV�-N9�nl0�[�}_t|��ws��ZQ\���'mu0j>/��H�.B*��[���@�s��N=kGp�+��.��i�"�#��֒ �a���iL4y/-A��N)����7�q�/��r��]C^DbGJHi�s�>�Qn^�@2/��#�F!ak�r�ڶM�1WԱ��Nb���Z3������X��~�$Ò�Ru0T��u�S圛\4t�:b���v�@��Si��|l5C����&Q�/��$"aG�
�ʼy	��u_� �hL@0M���l����8�,��F�W1
���X@��h������e�nzü�U��N�5 ��sq�F�!����� Syנ4f�0�[BT�ޢS��� �#Y���;m�P���=�[�.��e�Gʹ1�Y.���72��*��X�sZ��ŷ֕�wh�?s��������@&+R��Ky�h����Q�M�� �h2
dw;Qw?4)��p��( �)���\�Y$�o^�D�$s� �;_>��_Ŗ��S����w'_5�b�%�ǦA�<In�Ҫ]��O��0���Q�����XO��ɕ@����sL�5����!�х0��@^(J�����m��O�8dϪ&��P27�����т�1�n5�;.o�����l+y�ǃw��,P�}��i��)ReU	�l��I�[�ԇ�|F��{iuJU
3�T�W�r�M��P^�P�Y��}�@�4��
! E�`sO�%�m�]�E���P!:��z2�\�8�MM�J��U��[U�X�o�S�@��t�t���s�ᆏ/,���\�/O��{�7�sQ3����`�/-���e]��%�����8F�V��Y�}�(����y�絁�T[��L��ƫO��:����5v@��ӯ���HVЩ82��3A�y �]A8&���X�7��)�v�����u�%�3*N&��V_,C �����i7�o��싗��y�9 ţ=���~�,ٗ�	z����׫���j���J��Z����b�kY���?��Ejz�>8�T�e�֥����N����ߎ\��~�]�7��|��'�������*�s%�n�ysTOa]����6�pf�N=���zuuA�
��Տ7���yP���z� �3Js��w��0��ī�0'1Ba�����s�y�2�.��X_#"�܋0��ێCü��W�9���V6H샟��re�%:Ʋ6��% ���tZ;�RR�&˛���?e!�r.��|�W�bܝ�L��f�S�j�;�6.���͘	�р������JO�
���X+^��C~">��F�ȹZ%�M��J
���8q�Kb"�	���A��Y<a�Jt�I�e��6u#���k��0��S�7Y�A���'�t}�RJt���"H�/<>|mi^�=9�4���D����Y����W�:���F��g
�S�Ȩ2�f�խp�ډG���,�%HZ9ٱWb#P���~@�V[/�R�h8��G�)I��;�� �Bz������X #�X�`�}�hPB��$S� b�!�!Wx0]�����2ܜɥ��^������n!�L�D��%�J)S�<�}�L�� `%S����,����e8p���՛R{z�P�DК�0yu	�lE{�*��p�ɢF@�C�YD�G^�3դ3j1��+���"�m�I�\ ��_�f�-�ilOhRK�0��o�����P��	zB�R8��8ôy1���F$�g"��=�A
����,��k25Lonh;����o����jӗ�_>S���sDAz��K����=�e����S�p0�-�=^z]?ͣ�{k���	Ta���Z찈)`��WI����ܸ$5q͍��~E�:y���	�8�vJ<�l��l�,��}r;sV��vf��tV��BgUV,��]�a����8<	;6����i���)`��_�g.Н�0��]�Oc�K�o�5g�(�b���E�x�+�3FU��O ���t���l�4�E��c��Ĩ/��UȻ��������!��
(;w۴#6DH��SP䗴&C�ip�[0kc����"�6;���4�Ғ��r^.�y�F�M�k���<Ԓ7[�c�mpF�0^\@��y�Pn�pה�ɨ���� �%�?c���f��U)��	s�
��=��[H�X��S��m�+e�/�hu؜+�n�4���J`�c�Y�m.l�p���G��T?�)�����w��4��\)�Ci}�MX\��g���^���k>"P_I��2�>�M�dH�^��ˍ�d��:�
V?��EH�&i���f4X�l��B�,��B�9SF�h��L���Bkb.�ˡRq��_�.g�v����0NHP|�ڬ��Oi��%U˜O�/۫�WM��p����H��tC�'(ZV�ۢ�����vO��O�h���"�
�N�(�n�J������yg)���o��1@o�"X>�n�:aDJ�4W��i0)�ˇ�h�֫�;�h��+�(�!��푞ƖF�������v����j`�/d��>�%�E�eH�n=i�k���38��Wfp?p1�	�'l1�B �ۑ�U��[���"~�1���m�o�f�;�`���=>+�:���o��}�Y�ߺ�[��9�(�f���ԣM,󸳬���y RE�p���Uty��d�ki<O���j�shzM`|U�]y1e��ꏫّ�'�G� ?�	[�pZ1p��䀒���TڭQ�K��=�VW#�QN��=/2k��J.��@����T� ��Bsc�.��]�H;f�R���,Ó~`��f�����jT����{22�cYVH<<ڵ$��>� �����z������K�C]c;ſ��5i.~L�m���ђo"k�����%�����gu+D8r��-Tk�U�8����"��`(�G*��9̗�i6���N��>�\1���Vql�-�1k�yxa�
4���_D����!���LVV��G� .N��q���`vg^�����	b��\Q�a�n�JŴ�<��c��A�=ɰ��+��x���S������|�.z؆i�=įĉa,�m�Hh?��� G~|s|	���óϾY�?�E}��V�悍SvpT��#�x/E*�Ns�M�Fr���@{�h���	4�AQӎ��"ٽ�63��`���`���b�Ʋ��,��D��f�bG�]Q S�'5��ߤ�V�͛e��2�č��#)_�3�i�p��?��f]�\j�w���|��Ѝ��h�K�_ŨOG��8#]�58#�pB�a1y���vZ�dPy������[�ס�R��'c�j�M�%�`���(߇��k	�Z+`������t$~H������5ƌ�|�3-��aY=���f�����'�B�y�B���:n�U�ݮ���-���O�y��Q�?����߄����� �9\{w��J�^;�)Zwj ��r���X�mFv�d]�(�3�)������Pƣ|�EΗq�+�@�/G��M�����y֘Y�:�	�E��ֱ�O�0^ԃ<U�,��m����j������ѣaOK0CL�|d=���y.OӤ�X�dy���}&s�^L{1��T� �7���Xn�(Y����:(Ol��y oڂ7�4���,A}�ܔ]u=�EF�غ�_�T/p��s��������.pU�v�':���r���[]���'�?�?����d�^�0�2�h
�OЀl���?�{0ģIEo��a��i��,�o_��r�N�-�m�	�Iw�>��щ��D�@����,��{*�2�3p%���F����6�	a��m	�N��KU8�E̻�l���	����P��� .{f���偔ھ[ߓ�K�K���8e����y�\�7���%Hp���I�r�*���H����,Q�&���ER)��wҨ�㼤�~�I-V5%����R��e'@⹈�s�rZ��S�Ք+��l���[���Y��~�H�+�A���i��CE:�i�U06�6[�<�/q�'	>٬�C�`��P�{���`^��2����	��6���R��%r���:����yxQuX�%InX�-��GJ���-������$��*:I�	�{�ڂ��j$%`Iag0��b�%^��jMm��M���S��t��~��� 1�|�++�c-\�����xz�\�,*�Å���}>'�¬�\hZ<���j���b��p��T6Tp��G�쁘����@�!�z�B
�n�����]���N�yh<π-^�Ӹ��ָZ~�����x<\�qF~�.�������zrdg���Ж�p��aŬ}4jT��N!�}u�Cꩤ�8i2n�}��>o!�4�,���o۫p"�Z�D�8e�x���_K��ˇ<��y��OL��S;6���#���D�h$�9Z|�����w�X���$7b<�^�gF,���=�=n~љ�$����d�D�9�nQ���(X7rr�@y�5S���ZB����ɂi���6Ƨ�e��ws	��P���l���?S����!���0�g�D�p�L�N^P����HұO� �xx��Ix&o6�9��%4�ݭEv��:�̺ ���Ye&6������!~��W�3�x����HxN�3�;�$�����y��P�>�(��������L������� y��S@�(�k���&�g��Z�[�oւ��3-��FY4S���f���z.�Q�k���af�����0r=�w�&����n��SW�][j�Ln��b7�$��UK5<��fe�FfC�,]��o[��0�#��#0(��N����&B�� �Ȭ]`R�ʧ�5[o�[Aiѧ`������ÞQD���aOrFm.�<M�49���
K�D:���e��6z��-� �*e������t�x ���/���Ҋ4�����`�4���K:9�uq:\��_�����u���uK�� �F�S��E����B�v0k�.Uh��d�]n͎J�P��H�p�Jn�3�v�*d܄��zF�Y�mzQ���dV׳��$8n���}\^ey��5��GGa�ø��c���&�V[�k[��Rvڪղv�x1��Wð�uϭ&@��T�8>}Q`�g �P�����a+`BS̼�����p���c?��a��IZԞh�bKHZK,�\����i
�4{�ŐT��)�����)���|uzK��96�uz��P��^ �>�f@�܀���iȬH+X�"/iՔ'����ǘ���Q��W�uk�el'%���g��>
p��vŵ��X�2[Rߔ S@��<y��@�����Ά��IĽ��1U`;|  '�d��Gؖ�RN<����3����jVu����K��˯��ɑ�Tr�.r½Pr��t;�	~�F�|�l���	��L���o�c���"�J��Vj}��v��_�7�pc���x�2�o�����B?W�M���E�e�SA5|r��i1(�\�=\N^jÚ��5	k?�3�k6o�����؅f3j,�%ķ�y���4�е�zy���H[Q6�I�t˛����*�P��M=���u:��߱?���D_%=����ؑnHup��wD��_�2#]`OǮI�@x�1���!e��J�"+�u.b�%���Q��k�X�ˢ��PK�o���&��wU{�bBHܼ�b�]�,��"%whs�)`��'` ���L��ѥ��qV8e$hW��9.ˢ;��`�Ӵ?iF�Qay-�L���*��C@��71�if9X���m&�E��ٹ��U�6L��JW��m�D��tU�ZL�6������Id�EH!�c���oA�|�f�{� C�S#�7���R��x�K�#�s���&4}н�/#hx�����Aß'���+��9ʣ����EL�@V���_7�1�7� ��D�X�J�?dYXO�����T
]ų��~A��5�"�@3&w���!���MZZ=r�n����D����*F��� �Oe��.�{c�c�%�
�2	��~�/}��R]&S'1��FJ���kÆ8OT3�Boc�����%�/���ʑ�(ի�D��w�����X����^[�����$�;����zo/�+���:��׿�0o�7B��4l�rL�2�ś���4χg���p;������[z��U�X�gt� b��0�?��2�$N��p���;��,��%�����<���=W�OM�+�P�I��!�۪���vw78k3#�U8����ğ'�6��Z]�L�E�����B���-�5�����d��i�ϒ����cK��]��d�ej���o�_w*��w���0^��p�:�$����f��I�qjp�SY��-ll؟3���a��8�K�Da��_���Ġ�r�qi��	�����G*�@�T�=�����ٻ�2SÃԳ��YJ��膜�1"�}K�:-�*ۯ�����'�]�&ͅ����$4��t#g�YH-�Z� �'�rQ�P^�gْ�';Kݧz$5W.����L�̞�
�c����ZMZ� N���~��D�@s�,ؘ3���GjP���K=�f�J���0h�+F��r��jK�x��o\��d�EW�x���IWux��F[��!S&�)���=�|p����/Q�9]���]��� ���+j����L ��;���z���I��:P�:̗�U\��d�>=ڜte�g���0딜@�$�DJaf�w���ٰh��2A��,�E����ҵh��{��
��ʻ`���@�;���Wn1��9�s�˯\#߸�&��C��}�D�Z�"<��ɺ�*�g��е"�ҳ�O�.[�͗��҈	��z��y�Q8� N�aL�v��%��� ���{���pa���h{��y�%�O6K��#@��!��?2�<����1�&���۪hE�lٹK��	���.:˘�u#d��l�0/�P��R�M���L�F��
��f�d��+�*��*	��;���6q;�EP/tK��m�n�:�@����E�̾��O�̸�������TH
]ݙp@��ᗒ0FG�5穏��;{pѐXz|����|"���ć^d�j#\���P���*�����C�r�f�6�����!\d�}�ܗݜ��'y�P�]�5�a�J���N�HU+	L�������{~���s[6q`���ЖG�^	�E�%��{~;�.��^ j�"����5j6�SE��`���f�~׬*k�`�.%�P�wZ*6#�3��b~D�4�h�Z�����F����E�_���)c�(K���?�Ϗ�x�w V��q��U��0������'���#.�RJ��1?'X��T �3�yt�\��~!aW y]�.���R�������Q ��%�:��n7;���Ϣ��q�,Է������n�hO��f�R��XsF��єv�H������]�O��F0�=+5���F徘I"Ժ3�PS���x�EO�[n��/�,�{�||\^^��j?*���bvI�6xd�O���.���&�ç���"�:��-��$�E����Ѷ��4q%^�A������_����^�Ԍ�*�����i[�HC�OlB$��D��E+p�E�	��:ȷOz����g�ƫ�a:��GD#��sK�i���?d{y�`vP��O�C'fV��r�>?L�k2Je��b�ӊ���λ
"�Y������L��T���,Y�S��l��k&���������Ɓq�Qo���#�Y�����f�	)�T���fm\j��m�9��r�_SF�|]�}�4��g�6ڣ�rBL��Jb���&0�B��{腶���Q�N��Q��X�Gm�>N��v+d�6��_���!kf^wRA�=+�$�B�l�t�Ǡ�<����#`���PO��r�|��@!n���f�y�W	A��t�����q�ܙ��T�����A�K�Vv�H�|��鷌�-��w�h��8M�PеAc�����|b��.�bS�Kb�.k��q�9�Ku�MA!K��#W���5�I�H��zl|�S!J��G��9;�u$���q��}+q��=�KeŨ�V�䋒�a$�1�)~l�v���]6�
��ɪ|G��hH]��,6py��i�����I�8�R�& ��uw�L8�t|2�${���#��K��5Z���k�4��"d
%��|8A��}>�S�D���!4���\}1g�5,��|�@kc�Ed��	����ԙ@{
���k����/�Xq1�	ر�qVt����:�7���R��'����NaK��Aj{��E~�3�0;�D��9����:*���)='�	V��5t���u� ���9��P�I0�2�-�kd���#�|����Z��^�~%��� )L�����Z�Y�$���.��_R��{}6iZ�̧�
�bjȝ�ZL���	���;�I8�iѐ4)���t���E�!zs��wo�Y���;Zr���Zq^~���E�p�ĥd@$�&�����D��}i������\�@G�׉Κ���ĩ�>a���e��-��5d1�8j���
�E�U�{�/\f}�U��+g
=�y��j.�z�Y�b�f��9[��V���� E_J|�a�X����Z�X����[��������jT�ḛ[��ɾ��}NX�d��/Z{�!&)�����{��
Z�?��ˈd�}�6K���E1;�[0�&ڞ�������a�ŀ�mT��Wx{�.�ؿ�l���[; $l=4�$gҏ�oz��Mn2ք��B9�W8ҏ9}�Y�3qG��hVH.ݍi����?�4	͚�*!����ˎ0��p�3�M���w�76�ΪT�6w�Q�V�uSh��O|U��y�����B�Zkbs�&{�RLkVV�K����+[����������8h�+��y\��o��C�P��滰(�s��^H�C��\y[L������~X�(tx��e�Q��n�J|O���4���Jk��R[�}h�^}��s(L����10v��?�i��]��:�Z��O��W���E>�Z�Iw�9m,��{��QX�;w�+h��eī�C��j �ޢ=��ۺ�G��Υk��n��:��osR�о`OĳȻre�- Ü���Al=V2���)4�v�pJY�fʻ��/̦q�}b���� |O���?Rr���އ�
2xΙ��Ww������Vj�L �8]�׊4�����k�#q?:���i�1r$�rYS鑌��<Sb�L$ä����mR��Q��!���$�Ћ�K��v��;w�G���#�T�����S��a��fVQ5�ӧ�5�F�[��}��䫃#����m9�W�:���ū��]h�����5�1f@ߘ8� �����{�h��.��ϙ��i���
�c�(8�W|�N�@ ���+�C�}d�5��'c��[�D��p���f�<pa����F*3�od�^�k���,��������~S� ��D}1� �I%��z�Dc2y��F�o�F� ������p��-�O�%#UTCF���2��7�
���̸��q	���Jy?��c�b�;Ԓ㱌���U�y�<���-�����A��=�nM�:�b�$��I��G���Jun�wǎLCWu:��-���Q;�	�����Q�z���n�n�`#?H�����f�7X'%�(�s�/�S��������G2`aD�\�p!�R��&$�X�IP�Ya볒�3S.�u`ba�������1P>6�r��cs�P0�[��"���k��	p�4�3��{h�e�����;y;���(�SA���E�.uh��5���2���5����8$��Q3���" 7blr/&���<�.�#~ըt5_��Q"-�᭬zAgVZ!t�;O��1e�h*�r+�Υ<��6�y���1��W�uxa�����D������;߃��@� �O�n����hůC�,��D���=�&W}�C��ti�`�7r&\r���!�j�/E��qu%�_V��
prjG뫒ӱ�x���5�p��b��c#�C	��ũ�TEHṣ�\\R�����y��h_���Ffcuen]�S璿�-5q�p4�1�w�.��� �;s��A��<u[�r���R_듐�Q۬���a�jb��(Lq�'-kC�1��[�,�P_<�]��&�l���!��It�|��Y �OFъ��ʳH�gv(|fQ}쥹��o�~�;����^���!�4L����V�@����j�)�:��Xi�ǔUZjm�E��lS�߿�Ʊ?c�1�u�û8]]T����:�.Y*h� u���{�i�8�h����]�YA8j�$*�5{�ť/�Th�_sO7ܴF���y"lW,��W�1�-��%y/Ke�]����m+���-[3�
�M�� ;?����gb��6o�"�=j2l�~���R��Z"i�*]e�m��IR���񩛩�8M�TȖ�X��7x���.W��a���3`�B�И���ݽ���
3{�������k�e�Ūp�b4��-Uq@M���yG�%�K��5X%��W&i]2X�]�"�k�����^�Y7�%}�X�V����� �d�ƹ[�(ڍ�T�wD13q�34�������=	D��+6�\��B����޷��W
g�Y������C%S��4��J�T�JcpM����UP����C���B-<���xp���Ѷ���� �UAZPPR(ѿ��=��Z&&8ͻX�����A6凜mD,J��"��e�\x�<��i��d	�(�s/��U�G4ZcQTp�.��t�������'��DPx{�db�<���;%�N�x�>M��$���7��c��ι8v�����@|� ˂R��]Ip��7a:�Jīy���0y	�c?���[ń��[�׉��������c�6͂�Q>I�*�r�z��p#0�4e���7��:�g�GU�;C�i�PD'=]���5C�wf���h͊�@+K&�qc$� �r5.���J�<o�Ҹ��&�"�|}&Zv̨�2�
�PSF��`��P�Buc�.Ϭ���7e �"=?����@��0��!�0���k�5ͳM��d�ZY�!�؊�wգ�ΠSwKؾ�;��_�Ȥ��Ù�цL8;L��M�AawH��>�P�u�p� Ӆ8��|�L'���i��>r��;��^�9B�O��I}�,� l��D�(��V5���ݩ~Z�3�غ�S��(���p���v�I	��0����� ���Vx(�>Cr�G�Yi?��N\RvLO�| �>�z��eP`��C��9�%��'�\��,��E����ʲz��b�T�7t��/J�X_���?r8�K)h��$�у\�5�Zr�Od�fz�S?΄!(�S)�x0�����@�<��ҫ�e���ư"��J���w�(�Q3<.��l0�+�,��R��mr|�����S��n��i��z��	�2���M�����M%�FBl�r�֔�0?�����fb�S�\z��g7	[r�6��ݩL���c�T` SK�}���bi����g �p��S[3�Oôȟ[�V�׳�Y�JZZEf������Kf³^aP(���{���:S%(L�ow��GdX�v-&)��7��3H�z��R�O4
ٹe��g�����,K�b��!'�;8BDBMdm�La���#ȪrXV��0�}]�q\��v���Hb�nxk�����"C�h~Ù��n��r�ˬ��'A)],W��^���pPP�I12���^�G�ܴ'���)S��C�C��?�Nd#�v*���ڳݙFBa�<���&$Q�J��C�[��T�tj3�%��]�^�L�;[�4��탱� �R0?cD��`aa��M�Y6]T��M�>4�1|[)�� ��z���p-OB�Ϭ���6x���vC�\*��p�#���:��>��<�</��T�sy4�+`�땻a9;(��,a2�I�y��������{/�aD����7lR��Vf~�ǉ�2���"��u�޶��^"+" yi���s���'����e�DQ�ɮI���H�bU�B��L��_��a���Nb4jn��y�P�\��Ӗ�g�`��i�v��R�XԐ��c�p��n���"�\��[�����#:E��΂ǒx�9�3��V%��7��WԘ�ϗ��}t�%w5q�І���seB�PL���Rr��N^u��������-��x(,Ѡ�=���^�
+8��r�M�U�B5��⤪tik'����qJ�<Aƹ�����î]��h�A�ޖ<4+n3,|���=|�)9�.z�g����Уr⑅��.� 5�a�����Ӄ�>���_�����θp�u��X@�ÁĮ��f��^���F����0h�E�?��EC�r(� +��%u1 4ha���4e�(iI��k�������{�M��Uk|H"�`
����xE�R��!4 ��o��[���J�x$��l�՞z}P�/n��L-t�Hyj����G�4�~�t��!��9�"�a|vvO�U��dzl�7l1�y`��Fs��H�f��Me�'`��l�U���O2];�?�l�������$Yi?Z�*=����%9�J��~� �I�J�ab������Ψy��9��[7#��!�N��4��0���k(��I\�+o�gf�m�׏�t�P�꿟�{��ોϵyr?-#��íL�B��rS���H��r5F��D*��_�Q�@YA�森���*'��{��˲��DN�MJ��Ǳ��K�e4@|��a��7*��("˫��^�#�ۡʈ�$���2�;y�f�h;��+�SiWQt��9��AQ�>3�Ha��}�$��*���J�`{��b7�7z�RL�l�3�ߜ:��#P�u_��cw�h�(�E�����������i�����|$���5���d����ner?���is��|�&eUk
!d"8o�Y����@���K���B��̷E�x4���i��&�W�n[���ƚm� !U��'|gf�i�o�g�L�L4�.�s��E�D {��ɄB�=.���Xw-�L �x�;�����fML��S��l��*?�6x'��qJ�G-.� �����t��q%'�N�-'>Lip?���ʴ#fO�*$K�"h�)l����F0H�.|D�jϠc���	#�d� �m���Ie~1\�k�]��0P�W)���f�.2���ӱ6Ǔ�/	�����OH�S�	ǹ����?�i��	���������PJ��$���^PE��"�����M�����6�����t��IWI']3�wbJH��/���r�Jɔu
��<�jR��˸�vh-]R�%�9Bӣt��+�w�⢁ڬ͊�D+��H��ۛ��͆�"~�ȸ�5�m�L��o���Ν�lu�m������m��j������*
5]R+� ��T$�>C�S�ls9�o0P����3�V��7oD�|2�iJ�{F;�(�b�`�$r���GbUpo��d��$���SS���_��� R{�s����IԒ����H|���
/"+�V�sc(�3p�y�sz�U��ɱg�rI�Q{/��2e}
����r����Ʒnϙ����nax0��G���L��D_���I98%ܫI٩aU*��6S��	��8��
��dJ�l��jK�)������!&?�qWDwd�cDLĎ��l�C�?��,Rh$���u34�[Vb�Mj6eB0��^gݹ�&�!O�¥�&d��Up�4�op/(X�-�J�ă&2�����#&y�O��A.�E��Ԫ��M���3Ɉ`�hX���E]���w�k��;�{$9e���KK~���A+���6�F����I�KD��������v~��n�<%�.p]��.eQ&����;B�����.Ȳ��
ǘ�)�FkFջ)�j���[-��9�8�����
,|T=#����<���v�v6��%`ԧG�O�����As�t�[�@@GU�,��V!~1z�<�{�����rP�1��Ȗ�����j}�(^����)���R�5F�Wĉ��h�^4�8r!�~0��Ƚ%s��j�K�;��V����� �)#t��zu�'/���W@�E]~�>2U&-m��N�1��($��kڧ:����p+&�[+ر�����}�`	��O���Vٖ�d���Nk�B>,N��?
��w�m�Z�A�8a����+i��] ����.S[:�1�B��P�)�uwXL$3Z�ƍ:���β�bd�7���K_��{���X��������G�p��o^|��*���p�
J�=%��ؕ�ue!�Y�h��n�7uR�����sB���=B��l�T�D�?{i��4��S��
���:�!��O<E��ai�<�eC΋t,(�/Hn���4G�/s���ę4�{'�8\>fR
�n�0��C<f��뙧r��pv����{/1҆�b������-���9�{��1�^Qmg�lq3� W�DhP)�,�0�������9��i���_qjwY�eE��A4ef���i�~�@�U>yR~S�h�ϳ6�m������ӻv��]N �b3��x�<�F5RT�O>�^3���|���\I< ��Ӓ���ؿ�K��9�ZO!�.��տE�(\�W	���'jDp0�$���E+�.�H^�����Ȭ�'�kZx�Y f3��@N��~I��C��$���{%��P��K�+���}��u��Y0#a�Ҳ���ɒ@\����zݺU��-t�`��^��Ի�b�ŞJ�+�>k�Tc�eǡ���VfкZX�'j2�:f��rM��?H���~�TU����zn
����:���N���D[M��^^����DC�h rbs.M=��n�{å`X��-�s��P"򢭊	�g��$���c����(ت���K������=����0Һ?�tk_hp�$RdH���y%J��oۈ�'f��sC ��)A�u��C*1g���x<���xDU�/��Jx�w�~��@�wV���8+�`���t�����|�%�	�~��a�x����
�7���o?&00&.�ah���'3�8��\3�����=�5T�4�~@w������&7ə��'���� ���g��U!�̅d�� '���a����GR�,u�;�G�5�����|Zd	�q�^��B	�H�t�I#19n�t\��YP}=@4�T=v����3
%��H�q�D�,��Ƞl�+U�es�?�90M��ё��*��5��\�]4�����e�?1*6$/�\�}�{�Z�e���9uG ��ߙ��k{f�N�>��貿�,%iQӳ����r[رC?n��%d��ʰ��گ ��>[�Gu�4_aJ}���͈�^���C����Z��}]�WX��^�}<Bk���ͼ�2%�y� ��: p,�"0���p:�ɼ��q����_��#*�D�֭o��I���ԇw(��LM8�ZQ	�����v�	��GQA~u����n������RH%�O]���-Sm=��m����)��'�����x7λ:EV��g~�fV��	W|�]��vP3!�S�3_�]��ӢF����J�Q����{^P��ReJ��ca�o0`�&O�����5p+'�v5\Dޭ��T�8t3�����<j
z|��F��5e��.��%����/�M	�n+�n`���n |�m"�&}�k7�\�QC���g�$u2w~~��ogF�z:"��z_��d�!H�_΅��5�\�F���<�jXfH�_D^��5�O�+�J<I^O�~�gC�p^z+=�}�	�^-��+�T��7Ľ��#�/q��/�@�i��)�ڞ�����Դ>���Rk�D;\3q�/�eĸ��\��k�%5`K��W4��h�]㴇����j%��s,!/����s�&��CgX�8�\����.NF��S��9�����w�+&��}g�
eK�|�d�����b�;���:4,@�ja����i�X7�w�ɥ\M\D�m6Q�r�W%�q�Y:�"�d�^s�G�)v�f�Vþ���:���Q�M~�;�b`�K��Gzh%�,#��?D����kͧ2�t̂4�!1�Jع�
.��Sm�!>��}f��W�cww���G�
1�t���CD��@�L��A|����~����I:0Ty�m���ڷ'Uѫ�?�0��k�y;�$E���Xs�����,���l�Uxj�<I��G\"����]��Wc?Jp}�Q v�iD9���F8�,����;F�#�1�h\�;DJ;���2�����.�YP!�p̪�ͩq=t����^_u�+�#(-�B��TW�̶d߸��S�Y��;1�Xa����7?#���8#��tԾ��7�:��������!P�^U�W��MU�y3lp�� \rw�8�|��t b߸rA�;�����]�r���{�Yø�'�S䓏)�Dަ!�0ؤ�"m����*��������Q��f�﹟�M�z% ~ƽt�>�����k_j�5=Z��zp'���;�KM�g[�贝k��V��̓�����yI���O�E���};h~��$h��K&XM�Nj�Rÿ9 /z�f���Í�P����� �A<��~��o�14ñn�o�*?�3��g��(���"MӜ����;pyC!�<��h�k���$}���� m�8�~ׅ�w�A��ob�3�?�����hb2���S5�H�8��;K��#��G������
���|��F�	�/�\J���Ǜ�Ϻ.��˃(2j�+�Qvq?5�s�S'���	�8��/�T�kD���/�?&z���kگ]������oYڛ<�fX���z�-�M�eU�g�Bq�S]IH��ˠ2��%��75����W7{�����8w"�|��,��D�6��
� K�񗝾��Q�yt����ϙ�V��kiJ��렰`T֐Yޑ�-�)V��.��E�O�@�l@��a��ُ�;��5���x�݅���VNP��������q�@˔菙$��~����㷷iA���o�ˇ9�2��"*0Y+4���g���%�'�9�� ¢H&x�A�
<�.P��.7\���;� �5X��`.����u�-���3������`8�W{33u���k��dS��  ���ok�ԇ�d>��΂���L���p�?`�	��T3(m#x���u���e׉W���c֚Bn��;�Z�m|V6R*�/���5���>ե��ߜ��ߩ�f7v	��UTHl\�!ӝ
U�*��,���iҭ
4��8HY;,׸���N}4����t����x1���; y�=eU�����CC�<S_N��;Y�[~SL S3�LAɌ�X��F�	Kv��T�"�ů�;Mx#"��,�md>ʴl��5�w?�!��U��?=���tͩDk5z���,?!Y�ʴ���Rux]6
��2NHY�%���uX��}<R�}�#7$�`��'}�������#�T��Wo��,[��]�h�5'�Z����������rVD���d/�T�<y(_L���`��
���}8�cq?�L��s���T@���zZˍ /!\��������	fP���g��C!|���Kn@5M�@�����2kк�4,�i}�
�0�Q�Ŀr;�Q��`u,�#�`=&l�|^�e�ȒĤ58�H����};��V��=�,�Á�L�O"*�_O��~�%�����XR��'|��N�z�Γs���جn� -O��[44��VfvR^�xm}L�����_�ߣY3�����?��`��$#6�xS�j؝ߪ0b�����n%br+����a�ھ�H�o�5r�oˀ=;���Ҿ�NRv4/�ۇs� k�&?u;�e��Q��%�*��v���H��2����1tS�D�
�n<kv!s������&�{GH��r��j�JL���IZi'e�*FЈ��ʶ�4�쑼� �μ,w��2�׿�D0�-��M;F;��qc����PR���9۶��S�n���$�*5�дcjLHu�N�h�,"�OWz1̠͑��P�U��',��k�?|�ӾK䭺��UVrM��zx7�3��[��j�������!�]��lB�{,����e_~s���x����f�_��,d2!�ڪ��2s��1c�|�<���,��cC��H��@�dk��#�孠�Y�7=PE5�X�����̒܌�X|��g����óSa�2�e���;��X}YA#%7H�ڞ����D}C�94%�Q?��N��-�5u�a����$8��a`����G�@_f0ݪ���6-��扏�G��{��1��N=	���P���ǣ!�܄�l�na�%xj���a��X����-G��E���\g�E뱧(�͖Ld�~���+8K��=���g�&\eR_��Ok�[�Vbw���	��sd�-*��r��#e��NJϕ�=�8 �Jڊ?�q �aO�ey��څ�0'E�'�a/)<�a���]þ�b�%Eѩ���g�jg�
��8ЧC&�9~�_4��k7�d;m�|��='��c�YEk���To�	%�#��5a�����6�*��@�ͤj�i�@o��$���i-�� �)���A�!�G �4�iXp<m"
Y�3�s����|f�]]���"����]�h	���&R�S(u�焭Wk��d?������P�p��Ԝ��7�ύ���G���U�z���xyv�l��mt�V��B��������*j�#%�[�����o�p<�\!���j��S�&y!���/���$�W�2�t�(h�A�z�{�֗��h�-4/	��& ��?ܵ ���#jsSl���#�6�Q�_�t�俦V�Lwq���j�r�s�C.E��{��n�����bK�X���Α����v%\��Y�(��|w힜�������f�/Dw����A�%v�pwԅ���y|��=�e⎷Cy�  �+���,�,X��ؼ[�>�v�UGƯ�R/�T��)����6�?�˽����O��[)h��$�@�d4���.�EZ�Ã�f�$���K�D�<�k�W�o�n+��9��&�>6j����QM�؉�#����s��hZ�eإ��������I<?}xh�w@�i���>&����yen"T�k����)E\�۰��㈓�w��-��,j���,�XeC�V>���Fji��ܠF�	�J#ぁ�n��e�j8�Fa����w�^���F��r�D��M�/�����_QQ�]S���������B㮫�S���!�Py�*%{M\�	(5���8���)Ґ��tC�n�@�-�!њW6�Rtկ��9�k�,�A��Q��
�_�]���~=J���\l�,���ڐ�� ����a�DA�-�ʭ�Z���Y͔+D"�^�\;9�d@��~�]�+����T�MШ�3!���L�E`l�{�T,��I�}Uju��xF֝���:�ɥ$�W�|͟r�HZ�E	�����G��l�����eEѲNz'��0|��	!8 ���+@P���9��D8��^�x����lAY��XNa��Z�F�3�sY�Ж��Ι�f'�:����+Wވ�X���w����*�Nnn�,��_� dNV���P��S����Jj�AN�����
ZP���/V��h�[�:_Yp��ۦU6�!��qQ�H7��*������� Ck��G��i%(�P�Ul�V��)��D�|�u�?W�A�����Ƕy�قt$�~^O�1��?��{Oqa�j�� ""ߝ��c�6GA��Y.����$ً�|��H@M�Jn0�״�z�p�v��wV�B%��� Z�L~��F}�{X��?(�,*�(��:Oq�����xYt$"�Sv��x��= hr����E��$xf(���~^��U����DT���;�{���+)���ᬒ�7km����hԙ44���18��L��ޑ7魎6>��^��WR�7HG?���X�	a��a~A�`Al����d�5��zα?����.:����k�sۯ��7��]
�h����
�k�ב���yA����#DwwLk2����)�h泬a��$�z�qu��F��Y��������,Ѻ�_�_��R�5|P06ZQ�I�æ����ODM�#�ʹ=�Q���N~�
�����fTq�'.��#t�^J��ِ~�e�%Qn���	��	S�L)�� ��l��g+ˎ��0f��m��>����f�J�x�ަ@ƛb~ͼ�g�m_
i�0S��C��˄�\S�0^�������gQ�"�¸Og����H3��L�e7���Kv}�TY��@��ˍ]{S�.��[T���+Y�3lk���"p���C^U�y;��q�󎁓ï*uG�͙��DO�0�U�~��u�h�}�ϧZ��΃<TX����+�����G��{�Lr*�\�<`;��W�o�IC6$�4��amD"��A�����R�̔y����k��uB�Y9  �iش@��A� UFtS񧼪=)��c���en4��H$���Q��у�͝f1�#NO�e��mm
��R^#t�L��IUUu��ލ#QDT�je�^�ǂ�wd�~q��kmSWWߦ�MUós����qh���TPoHh%�X��[����2@�2�(DBt���A�(q�S����%LG]����W,�� q��Ioj�&���oθG�%�����"�c���<��FEu,���~wCra��f�u[��@�7P't���� m�K�>P�\2�s��w�q�{�鉻��r^|�=��w�z~it	B�Q���N���v�_Z�اc,.���1�ӫ����|�KTz'�@!�Ia���6"�˱d����H�i�.yu�1\����X����V��Y��s����u�&w�Q�@�y��;��A�B��M�J|�D�^meB7����ш�Ap=!�p7uTK�$B%��[n�^dP�)�]��D.>�]���bg���}���*�i�z��~��\�{q��:%��'mKXԎ#��.�3�$k��q �>:�}����:�Ξ�fB!1���%t_�?.a��E��{�h�"�<|�BF@��{Dw���[3V��91x��ɏXb��1=���3�.Խ<�����,��.�3�
q�Q��۬6W�^冀�5c��'��m9�I�ꭒd�>���<�����TWڴV
�c�v
���W�De����>��x'�� ��l�H8�R��5�h蹗��Q�p����bd�?���r������a��QV-3�;N裱$��VcC��Qjv?�۷�4Ć|��9F^���b�[�]�@^�{Wqx���u�(}HI�����ja�j�BJ���c9!v��8 T�}w=����q��P�k��ex)w�i�w�ΐH^����5�emI�*�"��\6�䄽ḅGI1A����"2(~�r��%=���?yx<�%�<�[�1S<���cyXD�W�7ٲx�5�nkfd5���cn����6�`p�N�l,���rI�q��h����R�F# ��vJ�( ���JB��B�5~�Ḙ^�B�B��(��>l�̄�;�vCq�z�`ty�����뭠�M�>D�RM�ꂫ��<̪�$�\������C������z��A��o6�{�7�p6ܦ��]qgB����kX�a�O��Pi;n5?���|�9I	�Fp�P��0kB�-�$ɺLxG��ۤ[�OnՃ\B�):���ą�n�ݘDw)������/�Ƕ�\�������׿��3-{������(?�������3׶�a�3�2Hud)i3J*ڛcQ�����Ob�v	����"�xx9����KAX[��7G栽��p��,X&�<��V�\pR`ܩ6��bJ��,�񧂈�f?��+��xA�0�2
�`Ȓ�\����l\�[t�=���8{nY� ���,�ܞ�t�WJWf۟?	�����QH_�.�~|Jg�E�����!\�EG������4g���mj����z�i��Ι�<�� P>�?$��&�4b�{�k����Z�԰¬j}G'I۱=��@�Ď"�R{~������}.��@�z�� �V��Bj����{Ƥ_�9%��"��}Q�������+�
��?)H�"�̅���u2x{Q�xhΗvJaԦTq�����q/l:A`�YΦ��҄%���)a�U�@���"�%n^�u�e�um�0yk��]��T����Z�#�
r���4�e�U@�h�R(�=��{v�����ԤQ������]��d]a/�C�<j&<sk9�<������ٰfW�+:a��møZ��7�z��-T�E+�\�c��=.�"�U�-�f1[U�BHoO���x�dJ�Y#<P����ڴ��J��l��Rm�����|��)��Պ���JK
��oPn�9޴DO�z�W�F�#}�(�O�9��Q������[wi�t8F*L����Wim�G�Vz�2�R뛙 ��.�,/e���Od�uw-�>�F&m�jA\��$,�����W���KuT�ʯ�XSg��*���O�$[�(�49i����SO������,R� �����d)��]]6�Bg�Һ�Y�NI�-�R��[��ۛ���Э	�cd�dUwnW#J�U0��Q��P א~fwG�Ҕ�B�7��G��S��G�gy�L�����M���<N�sx`R�J'񯅇&������	HHg��ܷ���o^�8�����s��4��:�Ec5�#I����{,j��06�lr��S�i�J�����.�韅6t�j�m�%	b��_��*�����"R�+�4���zT��G��`�~o�p�`R�ڋ˧n�[�K>�XΕ��D��	�YU$�Z��a|Ҹgj�a�>��n�	��� �XQ �WK�4���sF��ʮ$1}�*��m�{��h|.ot��s�:��G�
���ϪL�%`�c1��X
�����J�I�m[+w
&-3=�	xwd
!6��-4Q69O�,>�¹r�w#F*�� @TH��!'EtYm��8;��D����&)�n�jSl�E5��F�EG��p��Ύ�U��LAJ�6�Ф����2=��Mw?���ep�7S�V�o�|p��ARdwPn�G��G`� `³X� t$���ϼ�L%�Ȏ���9��*�����Ҽ,uD0����B=���-XO篚n�t�յ�1ZNB��.z��XBR�g<o�'Ô�:m��?b7�>#� �^?g��d߯�ӝ�p%J@K��o�9ܪX\˕B�e�r~(�AZ��#�J��
�ӮG�T�V��]��:=�T�ڮu�*�(���*Q���-c�ú'V��P�ֱ���V[DjN@ m�!�����Nc�"�o%C��P�-���%=(N���S�^�=SS��s���r�(yS)������?��r��hͧ�ۻ�� ��6P�^������!N<��6�{�p�"�[�<�7�g��B�٥��`	���,�)��D�/\�:(��c���Kf�ƹ���,�v œ�� �Hc ��˒����3���0� V��ћX�9l{�s�?�^���Fm�$��K	dBYGXNJU�C8*��.@)ފ~ֵ�6�Ի��n��fU� ��s�p���	-���|"�7�[ۃ76e5�� tt�r1�pN�e��N7lu���S�(p�r`Y�j���S4�& �<eu�>��*%��	:��.��$kI�8�Wb9�mM~&�G�V�1�9IYd7��2 �I���{�7j8��� J~���Ī�6�S?����)���J/ait^�v��\����t��x���z)��7��`.��lֱ�%޽Z��fs���VN͇ld�Ts{O<j7���ML�b��ʚ�p)��\܃�t:[�X`ǁ���O���l��_2���-5{���d�(a��.>�����/�m�?B� =��Zŀ��T��wc�{�K�j!�+"7��ݞk��%�sU�O�a%�u��q9Ķ��BC_P:�9Xnph���:*�tw/Y�?	� ��jM���ҍ�@��s���h��겤N׬����8n��z;O��PwvK�����=�kb�7tO�����Hi$��TJ�H�'��G��{�p��Wo>�!�������Z���'�<Y<X�ȸ`X�
��G4O�=�8�C���j�����"	W�F�|`u��5���NBA��\݂9M0����E�=�P�4�B���/HM��e����;��!#��*�A��L0�� *��ӛ*��K6��-���Bx���y�:5�0].>		޶��r�pă#���*��L�+�a���7�fJ�^�׻�t-�A&c5xyz�`h���B�˒��*5V�Ĕc�V~�͒�i�WA�7J������^ާE���(�
	�_�	�ػ��Bm�kҽ G~��{	to��VQdG�2_/����4q�Έ�r9��4�գ_����P%�C��r�?3�M.(+ �쓉я�S:ur�>�h@
ʖ!��(�����`R�䌟J����z��ǉ�<���C&Ȟ�q�����3ٱ�8�Xoz	O-��'�9����T�/(�c���J/�rkk
������-ZG=���OWnp��_�w��U���+���=�H��²�knz�w���G��g��q^RcKA�\=��.�����]��Z��i�1�/��Fv?�-p�
�2y}��� �ѵ��;���p�h��5���/NO��˒]�9(])5d���1Y�\��yBβ�05�?	|�����=�J�bU-�C�=M���e�+���h�I��������B�8�/W4�O�m�)��[P��٘>�q���Fױ����"�O<���o+ x$�D�sr�5��Ap�y� �ھï�'7� ��Ӝ\i�������@Q��Pֶ+�G5#0�IMlr/��E���p.:ܰy,רH���O�t�,���Y����E�K�\iD����*�Q	�MP�~k>����m�|��� r�2/�Pl�e^�A"���)�Щ.շېX�if}.����������o����e�@���o��a���jTq2��%T�"D�' �7$	��`�O �����Oi���I���?���H�w��������S,�*b����O
�ޱh��(G/���g&����P�gR�#�c�
������[e2"y� (O��dң�,OV?�q�6'�D�v����ۗ���K� �t�.S9,g���ɣT_w�3pZOW�]���E5]�e���*����*���:�'��cwW�}�!Eu�u� A��s;c����T����E%/��"����p]$�a�Ѷ�	u�j]����Xۏpg�j���Tg@�����I6�X's�`v�IaZ�J�<Gd�:M;7�Z*��D�X~��1+���������kC7�<�.�󩩼8�����J�~H�.,��m��Έ�^f���ܰ���"�j)��.������O�n�$.�A<���	'2�c��#��%���k��M>+�5w�5Q.Y�2+�I�{ ���Y�}G�(o,�5����/H3�;����7��M`�=��`8ʡ���F�Mu	s����D^ �����;�2��Tv7��2�R@4��&�?�YS���'�	�H*���d~�!EOٚae�Q`��@>&�ֶ��4F�}����C��EE���it[�5	~�m���טl�������5��szyP�p�sB�xݳC;�������0����ڞ��>�7� :� ��Lr��2I���Pٓ��Yͫ1�e�!���%��`�?�~5ҭNJ�</#��h׏nӿ��I���tW�n��6����6-0�6����9-�h�# ���Y�g�fG��R����eݾ��O����������
��7�4ah�+T�Z�9��	#��湮�# �hƯ�!m:�s�8����
�
��q_a^|)�@Δ��w�>��[�	�6���D %.�VW��C}�$�)@%��9��l�;{k!�D����f��FJW�����m.���U_�q\5����|f���3Z�v}���kl�F�~t��k�ɧ�ZN�C��G	Bh=������`O�+�D�.��u��Y8���ܧ�c�!�|藿�G�w�0"�^A�5)�ˤ=k������[٨
]G���iWC��'����&���`��ZH$��,���k�0q�wGY�T��*T�����!}C4բ�����&�������t��O�y��;�gA��%;ub���)�f�k2?�r蚨��݁o��3�Mg�=zq����⧤���7xXB�>W4u4��\� ޽U���
�-l��Jg]c�c��G[ ��]%E��ݰ��nW��nL�u�^���5gubNagӋ"�ۿ�������-
"s� ����
p��Ot����?���֭�j��w鏳˟��_OEC�����!���EI��ٷ������i��Q�E�ÊN���W��"��P-RY�SUb؀���CKsd��-~�yh�1� 6�;�/	wt�����&PH��l'�ٌ��K&��\Ӧm؈��w����/���C�0u9#H�H�paQ�rl�y�<_��
}��V���a��]���bX��~T��n�c
P����
�A-��%��!�"�RIڡ��q��d��4��{��]O~�P�d~6ƚ��k���D���ˊ&�A�6�X���o�^�h{���:o0���[�^�<�.���|�n\�W��mAa*�=�)u��AO�5� L�E)����r��J�{��q�g@y��*W�����;�f�-���<c�n`xgf~r.�M8���P�A�˰�]b�ZdyF?���۶�.=J��c�YN?�;���Owm�V�-xi����'�W��*���^T�ٸ�0���e��/�ӵD���ڨ���{"�!
!�+N����i9�~�I���PV�M9\��U��؂8ZL��H#ms(�"�("��gVĎ�9Lʛ�Zh�a+�W�~-�Z���������9@dj���+9�Ŕ���,�ݸ `*�:ٷ�����4�sQ�x�J�+�7��\  ]�$Bp��~\A�@:1����q	� ��?�`���{�C�4��޿��c7����p��,���l�bQ4���9���`������+n6��}SNL��#����)��
x��-E>�!l����ʇ��״�L��|C�Jƾ0��?e�0
Q�
A�C�G1�<9l6T��؎Fݓ��@1 �	=�?�����ZR�k�q�ՑQF5>[�3s�Bu�j�VȠ�L1T���d�Њ�~y�$���+�gI��钺D�M��S/���k�ߐ�\.z�3=����N��.��pB��禿$ws��@�U�:8B ���S�|&�z���1�� i�-t��WLd0DF�Q��ȿ6�Ŧő��n����o�}��IC<�Zw�8 6�"�m�i�/��N�K�x
��G��]J�OrH�� Gb0h�f-DE��������T�&QQpZ�Л��l���iK�jd�t��7�VE����K6Kf�P.���R�W������v�����jY�T"x��5:4 �bV��A���|Jԟ9��(� �F)�{k��6�B�����۵�ը&>ma�-��&wp��ؽ��-�G]K��?Z��Ӆ|�m�I�̙��Q����}|=G�E_#�tN+�ߚ�/��,#�/="�q|����M�dkX���	b�Ts#oRŨ�za��g���Q=��c�^�CѠ!�=��l���тr�2�ud1)��׷\k��+�8�>!"x�X�����/0��>��9۴�T|�	���~�q�_.T�6���c�e��Ӂ�03�������`.�J_X��Ɂ~�3�W|ج�A�Y�D��P��6׿��':�e��A�<�pډWG�}��.�1��jo���O��(16CY�����}���\	L�n�j�Gx�{)t�=#����\����a�B���g��4)�/�u&S�d�X!O�������>��(�����K�d잶�dI������&��ʅ|0�x(�Va*�2/cWܠ�������|��i�0�ކ+�0`x�<���8vL��Ɏ� ����E��e9r��ʾ��R��5_���6K��at����5~�%�kH���妈�����<��x.���X��A�G��;�֯l!M�T`�ÊkחX��T�����$��6;F8Y�m:=��"�Z� @ M�r��o�1���l�2�i�������lG+bD�=HI9!2���gIa���l�׆nD�=�@��D��5b�㗋��\Xg��E�	��KK���`�E� �f�8�� �e�fUw��D�q��CU+h�N�ߍ�a�u}�(���5|��/mzqR�@p��Yc�W4
���J>��c�|g�@�7:��#���ٰO�3���4��9�feKL�	;)��i�Fp5�^yQ?����U����x�R>7h$�rd�Y�y����s��r[��xpx)"n�rWy�Iy��5�.��]= �bw~�˕C%�9�f�>W����� �ɦ��}��z����!8�T���G���ݏ'��{`amL<��ې<�2�¼+�2k��s�!��6D\��O�U�)�@���-X+ӏ{��_�~���1<��
�>Y���B����ߏ;=���l�G���>s�Ĩ�8��a�*�e6�o]�"��%���s~K׹,n�h�5BE�t�U�+䣃䔖gL�|\  ~����u:��`�	VӘ���3�QM_��g�.���NP��Z����x��	�ĜC�H�B��#
�v����|�����P��x�0���1Jw��M6҇��{A<<��a���X�8���8��57�a78�d�%T�>[X&����w��-�a`�{O+$H��D��MĤ����=g�:Er
��"���	�]?2��M���0�O����u��� �ጫ�$s�X6L ��kg�3���2�ז#����F� �,ʅ��� ��1�x1�2��'���|N�rf�:D__�m��HrW� �'�C�y2����$�����7��<�.\�6�w�FQ�"���I���#fܹU���?��-��N9����O�?���/)׋$|Ԧ �Nm�?.O=f(�7�S���M�D���~ν3q�"憔���sje�k�<p�8��Vy�!�V�8�4���ƌn<��[�qk�"�R� ��9I��bdb(LЖ�~�;l	��OE�� 8�؍|��+�@CU��GV����.��[?s:^���Aы���v1|d����lV�i_;�9� ��Ù&�-��� lu����&�y�M�4�%2J���m���k�\[����#m��;������N�SQ�O��ʧ%s��6v�^n�կ�(��'=���{�4.{etK�!�G�TDG�浀�t5���gs�U�s���'5=��v{�$_�΢l�W*pS�����J�5C��
��4Z3n8�QcD��	�l18Y#QpҊJ����]�����~���?�2A�,�҃&y���b}y����p��1�"���M+?�(8I��-@v^_ zD�h%�*L����n➁_���o�V�_I��������h�p�+T�Ӯ"aL����5'���P3b�8�5wt�EF����IO�M;S��X�C�������3�[\&kʡ!���*�B�.�3��5=�/�+}�k�T��z�O)1��Ց�_j�Z��[���tK�z��*P+�JR5�<�*���^+-w��2�]t�v�8]�Q��x��4E%lnǜ�tOdj�	��7[���	�4�)�C�.��]�azw��߯��:"X����a�\ŕ��JQ\�7�h��Du�.��/F��n� =	8���m+�g�D�j�+?/�KX��O�[��S���!ٽp���;3v�X�RKV7�C��1
��f�@��G9��W��Y�	���^({P%SQ���wt-*�d�b��Szݫ�G��ák�k��8���`X�I(w�R�^J�����k�;
�8~-D�Y�>�v1�� "}���z.��_�$�.�V���U�w�l}��G����U�&����_R�˘F�!���	��03v�S(��u^��Э?���2ēJ���R�qQ���P|`&�ٴ��S��+5�.���U���O�:9c�T#��D �5E���(Qe���{Pϴs/��_���YL��a����zu��j\����|'�0��Ij�u�qm`�E�4�ٍ���P������I@�#>w^�}\S*Y�]����B�qǅws��c������o�9�{�'x.ws,牠n�����!�����x��3�fa9��%<�~ּ��)�o��w��X�?�\��1|�s�I�cDf�fb�	��^� .�xfǜ-=J~[��oVu�YE���D�����H�9~���r�N0��l[�N����L!?tm����C͗���k�Do���0]#?�`9.��x��FL�� �vKl���I���a��.�98&�� k��������{�x(��b&ޢx�"V�1��f+3W-������.�I#����h�	5[���L�Y�z�iCVi^�/��X�5���Jkz�EV��}�Ǎ���\�/��x��ƚrQA��^R'�oJ�	pĠ�p�m�ō�����[�"
�E�&��*d/�<�������Сxz}-�����e0���F����'��}EBW���%Ӕ�w���5���DT�����Q�ܘ����l^����Ve�g|�w�Cz�4�|��5l�	���*��"པ��Ws�G�}H��N�Og�C�T>�#_�z��?��8�@J�!,��e�t��h%��8D�Yfi����Y�l�h�$���E�I^3��	"���e��-�N��3�-���9��}iR�ϰSgp���n�����Ln;�~�}t������ ��\����D�&3)�"���c�_N�)W� �5ǳ�J����[?F��	Z���ң�X�@>x^�#;c���VwQ���
3"�D��m��pV��`�~l"��Y1��aUI!7���H�zt�V�2'9�XL���tJ�AW��WY�βғRbA֫MI�Y���xl
�����zX�#�!�s��2�^}��Ĳ�2v���*'� @h:N_��Pə�QR�rji�W.�6�ި ��0K�y2�in7�+�η@t!�w��L�2�ll����Lͪ4ݜ3u�K��ޛ�������)�ʪl;��7��n�!��xwe��m)�$��8V;���u+Xzn����,�M(�*��P0*�&�Tf-��Y��j��-o�Tƪ�H=v	[-4
!���ZTD�h���ء(�+K�NSX����q�Q�]��+ �ེ7݉y�&w�M���_"��G��]�Dc�bS�@�]:��E��f
DL���#��M"H{�1yR�	t4���*�:�56��`��E��/}��Ln�����lY�/�_{����u�`w����|��˺��	�f���\���:y <dl�[t�8�dY]��I�6�~:)�yj�co����2�F�!��gP�yB�C�T�#� 25:�w`�f�Qtod	� ��O�w�F�!�ʢ��6V-���4U���c�W�L��]�p�֜�.{�J4$�ÚMk�@BRI�01v�䍹�I�-p�ā��7��]� ?�k@�L���r����t�bk�d���|ߥX<yB�s7�����k�1/�k�F��>�3^�0݅-��t6��5�!��[�
I�ޑ��>�=݂���,j^�?��U"���kw%L���s�nn��i����]-�|ј-9�h�۬_Yi��P�OZ"���%�C��,5�jV������Q�۟�]R���bٌ�����?�l��ʴ���[7d��D.�(��e���;{��g��i���sI����"��0��ȓ����xj�qz�2�8��س�㛐� /e���:��@
߽�׭2d�,���q[�]�4m�z^�g֖�d�a�}��1і�'�S8Y��B�ʺr���A��MYBD�8�Fm�b#[d�4�#��H����l�p����d�bI���Ҽ����Z"�Wѳ	0ec���T�/��s{����z����ֈ%H)y@�T	�O���j7��3#���_e'9�Y� 97Q��5yYF�nM�s���}������h�
��`uN�C�F�&���^������D�B�3 �6$����9<�N�����lt�n�mdT
��X�c��$e���"ܬ���o��}T<|���e��j�/{�c�5��㥴C_��B��[97T��tQ�����{1?�哢�V�)�v�ے�5�����ݤ������#�@$����1�-�"��d|k� Y� �pu��_c�w;�?{�n?bief��rF���4"բ`�9�ͲR�*�p��c�DTq/Sp&������'������ڍ@6B+ӗ��1+�Kj-v\�sB�n�l"yc�6�L�ٶ�H�ɏ�����z2�)�'�5vRjj�4��ob��4u�m��-�5v��o $��N�(ԗ9�z�b(��
�������'�;�����$�P��6�Rh
S��z�7v���>��.�!�����4.�뛨�6��K$�f�^@Q�<��=�2����u�N6�A�y��Rܾ��x��ާ�Sr�<������5��rH���$��^��Zi���Oj�	���n�J���O�	��V zK\��zY`�4�Md���� ��nx�3,��rNtbE�Q�P�	�8�v��I�}^YZ�W���H��](�<H%��F�q�ǀ>Q|��(^ ��p�6��3X�d�S�pe��)���8� B ���W���X9��7�v!�`�vq�����~�ঐw��[}ͬ�ӂ�V�F�g������V���m���A�2�^I�qD�LS��K�d��;b��BfE����_�!|,���`�m��=�i3�Rl�ОG�X��o� S��r����Uܛ'��2Z$�޹0Ul<�3my]Xx ��o�!Tu�,Qg��B�F:)G&"��L��Km&w����>�F��4��N'�Q��LT�ye��x���SD豐���Lo�`� Q2x�����Eca�0qt`y+b�p1�ˍw�ߘ��NY���p���MဦȽ����k�0��#�ِ�s'%ă7�%ca��I���e�5������� K���\���V'0�!J��寔;0]8_<�i��,���J�Ȓ��# 6�a�g:���][9J����E�^#�IH6��6� 8�r�V���@����S+RL��l���CT��?U���~}I�@/�Br�:�b`�+�צ,&(�X㮾��U��#�ʬ���=�4��MԊ��T�X(����v�
u��]��`��Ë���dw��e��Ʃ�����z�"���vo�+�=@?oȎ4�$��#�	\���g�FT��
��uhgy����Z*{�û����݂�`��<}+s�YZ����8d|cCg�QaQ�
oz�n�%~�����?�><t߻�=�6�ۘ3�:�+��=�xtVOMO?���~D��BQ�;�i6���yl,^�Ҹ\�I�W-�p?L�k�,T�(��~φn�b��R_�����|�t½�١��%�IQ;z��LK�,KEB{��_�UL�Xno��c�>t�~�n��J���|����/��6�����&��r'���������L�>I�V�eo�j!?	�j��=0x�5��iF�-z)V� +C��K�_0S_
���l�xx	�G�.�����k����&�/J"�Aā��`�]Y/)o�&�6�W�B�$�~c�9�P�7v�o�}D�{#�S�8����M��\��	��d�k�,k`뫭S��I��jR%�2^�t�������Ggl��*8�� ch&�f��/}����A�ڎ�#c��P�� 9��Gu�V� �������R/>#ˉ=A�-�op�rӟ����L]� �T�r;C9-�q��t�{���[�'�q@	JT[���X��Sc�JYN��Is�dp��_sT/���~����ֽ ���I��"¥�������?���.���F�m�����.�4��F��B���V�Կ�| :������AQ�_���HzF�t�YJ2�Ȩ�;�^�r���~i���7�x`++Æ�iهn���GLuk-a`�T�X����/Z�]�(�ĝ�w��@Lb{�[�t�!�lؘH���4�|\��+�$�=�0rƕ����=@J���h����Ö�JKhG��{��R��O/�O�Ϡ��{k�؊��K����D�?qݶ%����7k�'a.Ĵ,�5�'g%N��sb3�H!6`�^���n�W�ʂ�4�&�?懱jر���.pcE������������q+! 䐗X��8�=��r�W�87`��� �x�d�sC�:���o>g�Q�������f�����	�P�R@U��3J!�aֹf�7�]�T
@G���W��)*#*�|A�+�r��3!�O�^�T*"�TWg[�Sן����!�1ڙ�����V"�X]��	�i��u^:�02`O�X���"�	F��� �G�6P�z�d�
`+n�?�-X�
�;����L�Q�Jİ���:�]��gNa�_�.�x��n;������ü�,��e(���<x+-\�o˟�u�;>��ߟ�yų�m��G��v�pk��<0f�K�W�2JYb.Wx���9�G�4+�3)'V�r��+�p�!�������7�K�^C���j@���Q=3�24e4�;��e���g
V�V cu��b��3�Ը�-�Kf�L_�f}7lbKU�����m�-�. �z�AI{iV@ٵ��ӄ.���a�4��~�%�V�[���ǅ0�[.="$�ܚ���I����c�:8�p�
���F7�Q�
MB�.6���.��J�]m�ִ�z�X�=��߳��Ctp-[��Js�nN/V�u�S$	_/���Щ�5��B�,6�
q��(���|�hD�"^g����p?��,�����	ՠ��mY�����v/�M�#�F�Y�������	J���KwO��\��FlH���$���0�f��H۵k�6S-.6cK8N�yШ�:��z�%a�4�0!���X��M5$�v%� �-Ē������L�1���V/E ��,�B�iS�
Y�ĄQ7�x�h�*o��p�#��%��p�}��M�$lbW��\X#�&[u�h"��N�����;u�x��4O�����l��4±�o�ՙ�����Ǌ|�(ȿ���s>�U����UJ�I�r��UV/�V��Z���F
ۙ�U+�uX+�R�C�R��?��+��s��ȍD�X���Z��rD$��|���ޥ����=�����������9K�9of�<Q�zR���s��w�d�.�����l>�
O�㳯�rf��6ݗ�S�����R]���M�W��~_�a�y�'��6T�>����C !m��N}6�ZY(Tϔl�,�
��
�<��Qׂ�Db�^�]4(L�M�r��*�Ȟ*�i��k�-�,��i&k�vi�c[>B�6T�����Ŗ��R���S�e}���~�о���ˁI_I�<5��xgiT�>˱����E�^g�|���8�r�ľ5q��q���쭧�1���I4G�2?�� tleGs��*��3��k���,�0�6-d�XR���X٘|�Q5N��m���l�ՎrdS��<̓��isN�G��t�X��m���c�bVU��O��#�:^x�iBU�{�ب�pR%����xmw5���K�Y��Dc���S`��]	�_���(�0�j(Ҽ�ݺ�g� O%��3�iF�OI�^��Z��v���Tf&�rw�ط����в���- o.�Ĕ��T�q�����է�Y�
�N����RAQ�ց��?���M�O���v�}�q*"3'l{�C| @�r�����`�G����gI���ȍ���i��.�融2���b�g�~�@�3�O*�/���k]�<M��v�eH9乊j� v�ٛ��yު�c�mi� AnƸ�P�wO�z[��>C��	uC�OG9���pZ�>X<`F[x��I��P:����>�6c���ǁ��YS=:7����	\rS~+������}��ڈC����Y߿-������J�9Z��_��6Ky�����zb������Yi�o�v<��z[c��J|�63;�o�:`l�WC_G�#;���JJp��[S���oYk�V�8�&.�hvVKC7`x��F-�s��J���J�q�1�?�C,������Ҏ���%ht�-.��N���׶Ç9�G���6;6��Yn�O:�^[@���6b���KCn�!�_��ݠ�ę�m��b��nʟa��m��o��/�l���kjމ�h� ��%{�2�_;\�q����, �&��%�^�|��Ѷ���\ϣ��zN�������V�~��=�fϹ!��l��CH-�L�D�qo��8X(��x�h�Q8����]*Ƽ"j�m�@�tpoY1ȉor����O �V	A�b��	Mb�ľ0Tl`�֠9K(�B»�����o���U{SO7�m �^[��w�v�rp��g�i�;�?ԀqId��G�h�Wf�>PH^n��s�P��*�4-"��W���Ru2�|����ه�
8�l��n�an\��bO������ʷ&�|BE���1@'��L��^��^����X�v�r��&]���\#��c�����N�է�~�)�*Q^_�<"w��d%����PT^�8�5��Q�x�1�]+�n��n5}�|�cR��odGK�!��S$�{�M�`_c�.p��{�Si5)E�;�����i+�2M�q)/���jF'q��f;^w~�8хϫǃ�����RL����,���S�3x(&��#��"�E�7";c��ݥ#�\X�:uN��i�kTB�K�Km�H���ŘO?j�(���u&F���,|z�4��zoX���[1-�� ��OƢy�6z9k����NY�F� F�����ث�����x�uqnIR�+<��1��t����G��I�"���dn�On�W����)���|x�{���Y~�H7��d�1�{y����Ǥۜ~O���t��o�"��oҕ*诮�̟��*a�TՐ�-�`��rBX�<C����𪱂�m���B�..��LNQ`����|�-nݰ�荒Y�y�#�����#���-�<$g50"-���YII�Y�{��DՃR�,y�$�GP<����^vQ�hd |rH�d��-L_z�dW�sŽˇ^ɢ�uQ-{T咱-��>fK�v�#�F#�1^�El[e��4�0�G]�����X���9��-Gu����Q6���Ʊ ;�ja2W$	�����A��J+Ȩ�<^/�U���c�L.�6��QJ@S����I�BZ<�m�3�4z�N��k'�_�~�-k Mt�������(4\2�qFp��O����4{�Ĭ���:bV^FcZw�n|_j]_�	�����Tz���<f%�xp��K�f	�`��b$0{T"t�_������Ϳ=+�
������]U xf�ᆄ���@bq�4���^�v��! �r�th���?A6�N�+�g֑,��3�r���3_����f�U��]�n�3�"�����թ_��y5�Z6��K>@�+#��F{��c��XTὗBi[q�%r�m/ ��|�����?)<ӊ�M�:S�z�J�(���u襚��8	�K#h�X+1�|���Eb���a9VqQ�"T���M����{��`1�"'��(��u���� �Fr���k�#z��H8����I�2Eh��+i�����6��V��w���V�~qL!+%U	�NF�va�Q�F�a��פ��f�"��p�=eR_�eQ��иT\���]�׿B��&�,v�`����4��jC� ;� W(�.�)\�1u[r��e���@P
r1�K)t߷�@����&�VO�H��R#1w�Rr��V�^��?����H�~t�B�J�N����xp
��YYI��^���nhq�צ�)q��ԏ�����������Ʒ�	�1�i)�P�Q
�kl�c5p��e�+�	Ɗ���>+/�?���fw��?��"�v���#��sSOy*~|I9�Y%��� 夙VkE��9[��PEd�Ms+�p��{X�b竞�wH��y��w��<feb͒]o�Ɨ�u�V���Ƴ���ǘ��l�Vy3�oC#w]��Y5Ŋk\T�7H��{I�:�`c��ۈ�c����>�Uόجu#�~���I��gZ�x��R�d���§��	�Rwb��nM��S�mB�v�49s��ы��(��&UV����s�t�m�eD:,ϜW_�a����z��,A�G?(�� 7�E�&��|��-�Y3���jJ��z������֟��1Mi����8riI�G @1O��b� �.�e���ҙ��kV����\���1���95�X��[UѰ�E�G��ɍ-^�Z�S��H��,(�8��o8�4V�H.��&�,���`�8�\}���ޗ�����dm*E�B���"�py.��0�HPiY�3�>�����@=MЎ��:9I���< ��W���e�3��S��R'�M<U�V��8��'��1cV�I��H���SFo;~�T�\�pg�w6�!N�3�v�T�
�r���
����"V��U�e��a	eE�oьH�T_�ᑍ0��^��x��;�g���ṟ�rh'���p�-q�^�h]�`��O�ip�w�Z�"������`��G܏-rd�d���·h���E������]�R����"@=2�|*��Ji�4_W�:�_�x���W�b�c�1Oz�Y��3��C����OV�\�<�O�f�qp��Pݛ:.�Sh#i��!��;/Wݟz
�ȡ:�%��ʲ�5�f�e���p�Sl��`�9��6�.
�h&Is�C�~�x�R5��P�I������v3������ň���e�{*n�w�pW-��eB��!(c�)o�N6����������{~�z�>KsN
,6����W�]�J��䪲ח�Wjux�^c��Z�˻�ԫ�#��R�&�X�N�F=f��}~�'Ni�C����{�!SB_;��Ӹ���5�����{C��=oe�	��ȨԵ� �7�c�:8z�.��nb���ח��hӠ���k�I��"ZvC�@�A W�{j
�Ĭ���W�f'G�L����<������:�"�l�-^������ca��V���ڥ�t;�n�쏧h���^��jKe��%��'��X��I4Y�a������N���k���n6C/T�/���Ϙ�y�����7�x$Fwᬾ������쩐���%
q{N��x򶫄+�{i	��|�w��9,�9T����|�Lp�a�k�u��B�SE'��h�wGf����F��3%�ĿK
�zBhfc{ꃙ����`ۯϵ�f��pT�|��{��zV}V���Ы��C����pS")4Oö�r��ruD`�D��m�z*s\e=<��)"7�6W��m9�I�kz�x�����8(1��m��`s����<�*�y5V:��W��?�QoO�$b��\�|��uE�H�ȼ.�����\�% ��e�(2�p�2�T�jݎ�x�W���ιs��Sf�3#��P���Ԙ�'G��W;��L 3*0&{�"�����	����}|�݃}b%�fii�G|�\���I�Z��A���v��\8i��G)��.0�C�IԖ�U�'	��.<��\{Ad�yev��9W�_>@�Y��t�M�icS����[e��X#�y^�3�S��TK�$:WY[,c�}�Ƨ9�ʮ�Hѱ�L%�2St_�ʡ�Ғ��_��{16Mc�� ��U<!aнoU��vߏkBa��|o%}_� �_q>�5\��~}
˹���{ �ܩ���o92 �ra�E���L�YTn��ef�l
���R-Kt$�Kܴ��ZP�)c�m[p:��R��e��ts5����� v�ߊ�� XP�?,{�r����XP�7�{=��o��srk�Ф�8P��,&vt�;�Q���)m(,CP�f���`"q:o�^�'s#{&1���`�6-�n��b��t�@y��_]��9����p��Ĉ�����O��Dl�]?�O���? 'I)p�=z���"��t<C"-�M�zD�&{�@\͆ы��u�gt�rk�%�
-��,!�g��>B�9Tg�,��&/���a�^�] ���/g�+�cG�tm�ē��>�님��q2��͟�>��V<�3�f�T�h���
-'1F{{f����jC��KRd��c(d�E�����(��xhv}6jYki'hL_��4�TW+�]Z)9$������\�M�$���C?�Ĳ`�'��g������d���"�'B.��#�5	��)�s�Բ��dk�;�\�5�0���Xo\pK��SG��)�>M$��CΖ0R�`ǃ9@��{ �l�-�Í���J��u-L�H������D����*;�ݍ%	*hT�g��#c#\ ���$��V-C8�.�"� ����K���(E˳�)����Cj
HZ9�s����K�J�[g�WuǎB�!$� nq���DEx:q����39��a�y> 0ڴsp�i�a�ڃ��Mh�U�Ŭ��+	v������-�l~l
Mni�:�&+c`n�5E�A�t�FH��|�#K{��٢�Dq���g3�&9*�0��
�^-��J �|u��%����g<V��ਸ�9��_�!��$)���Y���2uuf7֖8=P���URV_�����B��'Ͼ�]�SK2"�\�#��9@�q3�K�S(���C>��\�d��	Usn�ӼK�`#�F�\���"��f2�
{F�)�̸����`O#y�j���A���L�M7FT�������aD������O��f#	���:t?�ܪ�S`e珥��hXim��Td�]��O�Ǡ}��B�-�%�r蔠H�iԪi���嶄k�s���M�kV��[[���q?�?|	�-���+'ӐCh�.jK�5�Ky��޵���\��f���g��(��'���L���������v��уS"jgk������7�
m�[;Qp��ǇZhq�����;����:�����٬�ۗ����H��2'=��a��~�g�������I�wv�-�pȝ/:t�)d�^
+EP�A	�F����}o^H� ͨ���\���'f�9Ѳ����湼�]Cl9�vDNba�+i5��u<*�o��M�\#>�r��%"^	z+�$�S#�����z�9� ��yt�$�ցQk61��#�h����&�Y���0 ӟ�q�F�P�MA�2�����D�N�#
�+mٞaE%�������x�HTG2�k�8!'�$���IR�$n�4�y�M�o��� �~>�b.�5�e &��:a�T�bjq>)�~�N�����58I�jf�k��|[�X�U����R��H�ԉe�d��}o7#y��t�x�\:�y�&A>�A�X<͋_�Z�}�[�>�oQ���@źR_֯�Z�n��Y�&z����O��G�Gy):�U.��g������Kz-�4�|�-���!ρ[]�^x�6�9k^�^/��/!e��^�a�O��+�tʮ�no�-Ɇ.iq���徆�D�vm��z���6�qm�4�å9.=m�g�W�՟VYٔ��N�`��V�w�i�h�F�* (J.c�M=�w%yQQ@�>I��r����fނ�pXH�.;��b���I�R�y\{�6&��A�eqF��xe@噒�(�?@P[_��r�C�k#�G숏�%���rn�5샊��Ҏ�U���ݫg��&�S�s�����:#{��*{=�Z��U�񂡂�Sn&7tdD�̛�ළD1��]��H����S��R
;Л\!�c������j��w�!��[V�V�y1���2���n0B2�c��/��l��C��d��l�n�'�Mo�F����5�3�q9��(��ڶ�-�1�aezSti��m���Mت�R�I'�j� ��N��F��FJ�]4�jV�ٰH(+2���(-��v&��UG|��G�\����1[tA]�C&�s]���J�Roq��Q�Ty]�3H�]�BD��HK�n��v{i�a�W7*���U�X�*]�τ[�Z����N�:��ؒ�1D���
�V�7M��F2J�i���<�̀���B��&��HT��E�Lh��ڰ`E����JK��Y`�}�<L��i���ndq�$���⢑�g[�� ��R�J.������[[TXѻ���$��JCa�b�g����mƵp�b/dTǽcӠQlY�Q6 )�~�m-Y�ʨ�h�M��1��7�*�L���;j
g�	2c�w��^���N�L.�ج���5�V��� 2� ^/������Cl�4Y�.Q
��j ���!��o��YHX��ȍ�����Ǭ����{F�9wX����M˷$��avP�T�1/_�3l�pA&��X,�@�i��=56u����y��e��95D{8υ��Z���HN�Y=�pە�[H?XႷݧ������%>��^���hS�>�T0��~ew���[4��A�D�|z�#��	��c�~��ی�@�ݙ�r)�ɿ�2��B���C�<�;�ɯ�i1�sB�������٢6[[*��;��+k�I�/�h��@��%O���h���c�|�mQN�݀��[>ߵO�a���3Q���У��K-X���L��v��W4��7�.Nd͝��U��3�"����VUscX��NO��F���e�X]&zA%7�����E��o=�ٳD���6� ��~�*�^!:Ϗ��b �ҽ�#\=�>&��` �!S��ʆ�Tyv���S��+��F3۸�
q�qQ'l A�1� o�`���O�E�p�����U��f(�M�����WѪK��.�1]���\�3�B��k�g�*,��	�O��H�p��rH�q>�8V���MA��ø���Jp��3���-��J�K�;֊�a����0�Q�X��߽E��x�c��"t��+ )�*"	�����S��_~�-�N;P�T�1��Ȱ��P�g�����W9BMnR:��ă�(I%�i0!}�HxʡP��+��]ߟ�)�¥���ԁp�W�s���! v�N�.8D�L�U�`{�bݑ:��$X��na�Y=EF�u��t�><�������w��:l<�w�M�f��2+�Y����(��e��oL�$�bF��O�\����+�݈%�cβ��&5+�E�(F��c�`6�qM�􀁦�+.�^N���]���$V��-�wG>fI�Oj��8%�ݬN�pQ�;_W�>��q����m�X%�]ߴ��Vn�v�fl鲮s[U:�v�,�g�?`t�<M��H�UzHs3	r}	��L��Č�*�cV�L�h����hf}βѺe3�g����H�+��b 7�Σxʋ�'[��p5MT��KH���(O1�[��
�~���c�f3��ׂ�"4��~��_��t��֙�.}��Ip$�)lEp�Mt��JB[}ܙ�0LY�L�ʡ���
kz�1��|%C�%β�?Z�!�A�����u���q���u�e�dFK�#=��P��BU*0���2���8�hGnGh�"��0����|V�݃���ud�ϊj�"2dڙ܉PO��R��I&U�!��h�QH��mWn��q"L�����ןZ��t�6�D�u�ȼbw�s	A�TW �wJn�%�{��w�86�~7j�*�ӑdo�ޚ =�WFG�܎�zs"�.Ez�C�3����V\���Q�J�tI�0X���xbmd�ܪd}�(��9o�*�9�r�a��_7%64U�̴9��S��1�~���1�
v�~)�p��c�s��gEJ�sT^$+���_��=��s��}�>�&{��'e��9��N�U�c��}tM56o�E�5rq�J����1���X������M*G�h,�o��#)m�����wl�F�QR}k��Γn~�|��w�������hB,�l�i�*`���o3��|�+�B����$7��b���ΒO���<��yF �\�ce:<�0���}����>eSc�J2����5���c\�VWh�_�|�P'����M���
�����c<]��b�2ҥ4 4��WM�F!�SC[��b�����m�7b��c�5�����5~R���h!{��Z��_R?u���|�*��,>qQ�*ͦ5N2qʆ}����j�k�2��*]�(�&��d�@녁y<�=����G���I�!?B�H&��c��Qy�O����3m(9�=U|�@��YF�%�ɯ>��V��b����CČ����e�m���-}�W�������.�qF}:磖���b�+��q�\��U�Dm��* &��,)�]eE]�{�G����.�0��P��Q�M����S�>F2�aj��I!������x�!6ޯ��2�{b��l���޸|��r{$���b	i������:\��������*�է����h
TLn+����!��Q�Y������Q�o##������rf�A��{Ќ��=�x�*��!7�{%�ID���·5�p�����5�2�A<n� C*B�Z��I��7�D�-A�I���\"���i�fn�OW,� |:����\���xf`����#,�k����r��v�v|c���%i�CY�!�Z��6�i3I�Lna�;����1�#dc�Y��LEP�߅j�j�x쥬y"j���mx�ңVmfPK	�����  ��?��	���q�94?v�����_����$?�q!�p�G쏭a�����3Ю
�5g��u�g�ݶ����f	ٶ$3>ۿ*��9�6�W�x�ko)f�d��H�r�L<ě�	f�c톸�i-�����M�6����Z�����Gn~�p��B�Nf�G�V>f=혥o��x�P�fe�AFǄ�io��'��Ĺa�i��9d;U\�^Z���t������("����08B{+���P��O��]�V���>�qX\H���	xw��2��_����@�Mi�2�.���Ox���=��]P��7b-�^>y+�$��t�Jڊw>h���(H�@�dk�a��[oY�4z�JT���2�w����-7���]���׌l}머�6(`��%N8��sp�.��?�Rp
E�Fz�� �(�����y�MW���|����C�k@��q�hm�'Wg��
)u������
%|�I�	�Q&�!Ө��]��b�+�)	�I'��[��f��i���E�w�xu�8U 
�[L�۪�L�,���@��;1�K�-�ñ&`=���:�K0�dhN��z[ɸ�n��l�S$σ�q��㪣���<���^�������Į�gA�'�9�پ���`�HL0G2��#����(m\�&9ʌ��bz>T��ݓj���HC�F�F2*f������VPW�!<g���v����U!���[���1��nc�
8W���F_����ޢzf��Δ�KP���9�Qr3��=_U%-�5wK&�ж��!� �(x��������+�6	d ��%��οC���[�����ԡ��+#o���=I�,J����� :���x��d<\NJ���ZKE��Z��C�M�e9gv����&^�[ޙ=g��HN�0�����]�[3��A����鱝ﵑAGDj��~.a�c�������γ2(;t�D���_6u�4.s�b����0ɯ*믿Ð,2�9V��zm���Z��Jl�={�!��1�;~}|�v��_�2����K?~��
X�ȋ[�9�V�rI�0�7��>�z#x�����0�5{�ST�| 5�6#�gTa��gY����\7�l2Lѹ�0���9FI>0�1Zh)ܘ4f����97=7�a�*	&]kB@(�3ʐ�+B�x�����)�b ���	$�F����$�#��-V
3�e��$/�6@��髃�����"m��G""5�'�@�ا:��r�A�vNj����Qék�	P���ٗ��<�O��$�z`����]3�z�`��hC�����,i@��	�v���]�A�r�}/e��3XŊ�@��EѤ[y��w�2-./��v9q?��k_ս&�P�\1Wg��`�>^[1�A���e2�4��Ɓ�b{ �f�x���=$�L��R�#��j7���p �((��\���>d���PT��w���{7�m�Ʋ�w��_n@Q!��MX"�������n�Z�j�,��ۣ����w�Õ��	�s�~Sbo��~d�l'T���N�
DC�Q��?!�����
H�+��M���[�Jk����'NV���xp#G����𑇈�
�KU�"\Үh���0[�14���_v��o�>�#�F��q$#eվ�N#V�mQ�����tS�V�3<?�8;O)��u�
e}ȏ-����	Evs7Zw���C�#�{�o+���C|UB���m?�* Ri�ZH���ގc�P��u�o�Q�hJ���tMr�}�$��	��=|��t٤�1Px��n�;����{�VI�2q�m-����]��}D@ ���t3���vn�g��?�]
Ёn�A����~��p1�}�Iu�5�Ap��/�w>P?�Vٝ�F<���UF.O�&���YP�O���BS��� V�{O���/�6z٨��n��&zK�e�b[do�����p�Pe���J�~ж�S�މԆ��86��1&����ϰ2��Y1���k�E�T���ϰ�	��h?,�G*.C���W
��Vk���b{ �5M�/W�}��[�Ԣ�A���jq�_IG�u�3 ���I�Mưx�ʳ�ڛ���A��)4�5��1j0}�ϰ[�,�����:Cϻ>״͗e�wx���A�P���N߸S8�Q�' O`j~�O[�ǆ�+�<V*���k�?�tEM'"��Enɡ^��ƾ��K�Ӎ�2�o�	E{F�Ȧ��AC��7" 8;�?����|tf�5H����F)��r�"Ѱ�ޏ
е,�=�_ƝQ&��¥5^�Gƚ��&�:��r��vi8�s�9����}
z���n�{�аs-�lzvÂ����	I�O����!u0���20o�*�6z6xm��D�DZO����G����9n|�l�U7�|�~�7o%����=K;���5�� �6o�-* ;&(FDtǚ���,������|�$M��WcO@����k%I�\���jB ���\�߳g�x��T�O򈪢&�X0^S_B��&�H���qqT�xJ�a{wV�Z�̬̎9$F��QU�Ķ���%S:$J�8�"���X���o�
Eh{H�k����ip�폾�o(�`����V r�}@�����Ӻ�	f�1��y�����a(( q�{d����3	�`v�!��.${��^(��
M"��2@�]�[��b?�~nnk5<r7X���Al���_�q�H��6oC�<]7"گ� ٵqA�}=�6ӄ7��˗$���H�\� Q����� Wz�ت��W�U�©Pi�NP����[��T�)��VG�Ρ��S�X���j��R�A.��}f�y�)�Ǜ�%X�Q��ESGH��Nm�᧣�8�ze&DK����M�	R����U��e}�H�g?
�.NDcղf�NG�fF���/���1�~Sp6�K�Pk�9���t��rd���L�������{�Xm��{�"�8��;l�%�tdy谗����!'�jCexK{�n��eR��ad	�J�o�vXK�,�ӊ�Y���K)G��=E&���r%���/��(�B��ϯ����0!��G��H��|���Z"k�02���>�
9{8-�Ik�D��ǯKe餓��o����xI�(ȟDv��f@L�oV��@T�
J� 9ȯ[�2��.�-���u��uZg��g�em��f��|�V͹aD&�ӕ���9�4��痄Ql}��b�]�3�����ʹ��6�O���Q�-�t�ݷ�7'L��5��5��\�H�p�Iw�୑B8�Q��eFI���]�9��������Y��BV@+��v�{�����BF9�oZP�����P��;Hs��S��D�Q�	����R/h�o�\g!c0z�R�¼�1�{�ݬ����l�)h�I6���_�r�"�I�	A�,b���],,��ɯ;����wO�C�:�`��-���s;;Q�C�mO"�yvi�Y��)٬�����=�$C98"G=f�}v��h��a����a�V��Xqy^�x�2�� BZ����S��wH@"�pI�6����҈��1�At(㖐��Nq⼾"�1x�jR}`���Y�g]�ޝ�o��!�e�N���unw_qW���ب��x�nН��Ik8n`��z=2�z����c��B\ٍ9�
�]�"� n�:��qm��p����:J���=H_[�3��H�{/�
�<�c��������h�����7e�H\e�5w_Ms�~l��_�����d O?0�l>8�����Ve*ۜJ��c!�{xo5n�y��C�sFc���l�(�O�"HBC;��?v,mɔ��葉����n�,��[#Nm����ݸ��8�J�ܡ}�WGl��)��E݈�\9Q�M���y�7fp��X��2u�33j|i�L�8�U1�d�b4Ҙ����^]RO=��?RᳳhCv�M;ɀ�����n�3���7���
Fߌ�JK�Oу��j�X�iѹ���Z�~��2����b�IPST�]|f��+`ZYw���MF� ǥE�
,���ɱңR��N��VC�[P'NV˘)|f�����x�d���B1�]�k��#����v���!D�$|W�`�p�O
��e�@N����!�G����5���^����}�d}�.\8I^��|Y�p��Vs�eL�h�"t���oK����������^U��m(5Q��YW ��Y��CR���� Xڷ�V��7�Um��H���n��c���Z�Mv4'�Y�X�6����t�:h�&���\���iy1
�nqѱ/�wܸ�o�D���/��{�6��FL��~�]��m;��_�xQ�:on��Ii7R�^]��ɢ೶x�m��Wأ�H�!Z�#�8����韃1���(Qq�(F����3�GM��N���%���e��$-�ʊ'�}�)i��`��>��Ք�"�<����D���v%�l�Ѡ�Z�*n�W.Co4|������0����X���� 9(��M]��"
��W�|s��\�U1&���;]��$k��NE�~��z3�nN;G����M�C�	��#Б"~��
�^�4������sH�FۖB��@�Y�f���9�ۮAb���:Ӱ�wOQ
2�G�o�U��M	m�U7%x���XDu�s���l�fDY���$������d��%1ݜ���C����J�-��2� �?r52���?�	*����Ds/cw�u(|�}ٲ?Q�夰~��&���/� [ŶZ�At�Iz�Ϸ�,t�h3��V$��7����Fb�="��i��P} .K�jAk����6�I��qv�e�a���'�7K�����`F�H�d��f��,S��ߍM�4�[�<���k�l�~�Ѯ:�<,��*��Ŋ!c��[�����R�j�D�*Z<]�ɖ;�"���@,:	���x�����Z4j+ֱ��ʚQ�3������i����o�C�%��t� �'ө����]�m�8��1N�$a���X��AD7_r)�}� �+!�I���3yܰgڝ��9Na-|��������UM�=$]�x�f�7mě_��X����9>��
��ٵ`l�����]TgJpl5���Y1O��F#-�f{(j���HI�	���?q�����$k�L^ zl�u��|ev��M��<z�����-	�n��!Q��N.��m�H���Q � ��:�HVa��)�<ߣ��=_L5���O�j4k|���9.�M�3�cUE �.u����>���]����0;sj_g�4���-�W���o�	9wc-J9�[�%���t��oU���V"�yj�#����fvx���=��.l��ӎ//�i��Y�W�9��6���7�u��_���h#`$SA���W�A���lb�pΜڪ)gO) ��U�ǃ���Hm�s��H:_i�Ι��ת��bZ�I_�#J�ۓ^b�:?ͯ���~G�@�wo��oL8{@��5E�
�K+�6Nu�'�8�q4^W��z�m��Ӛ[@w֫V��$	P-�xi�#��YyN)\�@bԕs��j�H(��b�н�F�wq��SΑ6�=Pt ���c��-A���Y�+�3�y �5�2p�S��V�_@u�8�u<�YJG��
sI>M�Ӥ��������8�C�/��n�E����H圥�o��PI�Ad� ?��S����.�/or9����/�5v�kFpCyVK���,�B;D�t"��d�S��];�Ӡ�(�C����~�.�����a�o��d�j�&�Ƈ�4#���h�n��L��?���,P��o�+ݲ�	לd7v��6�_P�/���"��^'�d�s���D /��=�����q�Y%�FX���|��b/`�m���(<���GA2.�|�t�2��F3�6���[4�g�n�s�o�K��^����$b\�¾��=��d�I�5�e��l��j�t�jEl5��.(2=�����鮣�,���\�_���<�ߥ�p�V�!�kN�ᄛ��[:���b�zkz�໴W�
)�͈L��;��<KT;�)�O�'�>�ѻgW%�L�	�}�'0�ʸ�-�c���\��ŝ�Dȯ���?������~�'O�y�d��8i����.:����4�m(���y2)���̦ ��A�VHqU)w�n������S+��#�h7�Bt�BW=�H�t_�����y�F��H(�*,�۩��&s��I������1�%Ӛ^���1L�,�@��N��A #�����������5K�g����t��7��a��ԅ���DNk �?Y�S�SaN)q�@\`�c�Bc��_�D�k�!�&;zל�`���9�S9�ɢ��޳�ICs�jX��]�iҟ5��+Yi���!�JnF��M�&p��%6ҥ�'v�M�Ƈ���<��={�LN.�cU��{�ڋڜ�e#isZ��Dc��S`n{V����Z�I&gjx�xG|-L���
ŏa[��N'��k�BHz��� ����p���T�<�-���T�%u!a�x˴� ���菡0�UJ�VanW<�X�+�cj�4�l�n�i�.e7��S�|$�����P�[%��#����֐� �E�'�糊 eu`V���~��5#���L�:����@4i��X�����oN�\��g��<��d�`�@�𒕷2#Ю���;c΢�{��k@�2�NVH#�C�����Ó�����!�B���޲�R�ie�(��Q#���\Z�7B�g��/�J ����a�ʵ̭�����<%l�h]��}�\�
72�X�DsX�S(��+�:����Y�7�G�vQ9ӫ�Р��n1��}�S R�TS����~d��,�(�$�����1�Pb�tx�WTC��KQ�lF��&��ԁ�Χ��/͇妠!rP���+މ��DC��4�Զ!/p�o���r���?K;M�2��R���т?"g���7�!��}S=��8ix>�"�Q�м����lE7Z97��6ƾ�� /ث�q1 J����љ�S SU7�J�аdM\�(>�c�#���oP�Y�Lx�lpMm�n��d�`@�R��*�oΰI�3$�	�_��H-��E>,#��T�f�I�2��vМ<n�:w����g`�1��F�e*���֯��-��Ma��C��s��t�˛$ko�62.�Z�X`e�1���3�j�C��8\�%���V�]��'�3�!^9P���P'>ɍ��Ғ͡��χ;����W��+�)i�f����t������D9ә������U��s��j�a���b���L�=ŏi^�'Յ�:d���ch��Q8�!c>�j�+��)�L�y��^ۯ�a"��fe�w��L~���]@�;YDd�#U��6�I�B�������|�a	[LM�=S5��^�hC�j�.Dm��y�>Jo�Vό�Hn%�>�)`Y'��~�k,�c��$�<�$�`p���=�QbxP�h��:����+߉;�9,�ur�y���_���سɖ/];��0��u�J�1�����~g��R����"�|�7�mYv�ť^`{�������YD� yp�#����w�"�Y�3���%m���C��U�Ut�-���f���Ǖ�{ZZZ�v'>�Z)���,��1)���̈́��
U���H���{a(�W��OA	����K�˜8�0��:��^u���>Z0�:�K����^}nź�NVE���P8k��|4J�1��ïW[���#��D�~У�]�<�n@'�ѐ�M�(O>���N$��Qv�|�
b����4J�Sl�>6���U!I��V���� I�0��-�j���LiR���B�����R	�;;O�i�Y��b��syk"D+P=[K���>/'��{ͳq]=�f�� ����M���j\gOeO[���m3�<J���� ���R���n~�g�����Tb��'J���C︡Ka��[���.uЏq�߯b��N�-�W�����~�Pk�¾���{7��*B����|�e��]M��m��s�@��1��ލ��l���k�;]������{�R��9��=�Zf.�����t��Ẫ�`0����-����{\NO���
��gx���;K��`P��M]Q�v��7Ƃ��l�+�)�'As�WqH��'O/���=6�I��V^mCx{v��#*���P����-Jm����	��]��A�T��?pE�w,�����k|~���R!Eo_D���AR�~�X�saVP���7j���l�e�N������!��s�%�.�|y˘�?D�NC�/ۂ�X�moG6	n݀C5#Ʊ4++��Hܡ��H��������۰.���r���㒳�r��w�#GԪN�����s��V	��A:&����a�ɛK:S��������0R)��PXz����I	(�9~
�4�r���>=�k����ZUH�,v�l�Gj��?7��2�C�5Dq�I�:)�	
�J���ǝ�b5X�3��!��ZeH��
�;�Rk��^��cst̊�@���v@Wf�^����S+�>�8�^^���7�3��!X��Yt�4GNo��Pi���<��,�r*��;a��/�����?-�N�������*�v)f	8(nQQ���t�sl!ga:F!�
��}������*,6�a@�f�ȸ�t&� ��Mc@��4��F���m����)���]�f]��T�Yvo���(}c=��7{��Z����C�e�Y����'˩�~}�r~�����vp�}L-�Z �M"|�v���bz������p�:��~&�/?��h�k�����8�Qu���e%�F��x�!c�FF���_�}�׀B@@����xR3��G>���n�fx���s��c�;y���`!�Y�d�em��7��Z=r�A�N�9![����4<�}���tQ+����7|Q��n5+8�O�{[�d���D���C3�<u��2l�~���lj���Bw/���@�~�=���x�\�RU�����yX�XjT�,�<��UY�ek
�F�H��9��զ�(F���g���q�c8w�-�;�kR����BE@��cq�px4	�uc Z����]5"��7��3�ƀ�n(Uk��r�>�n"��"4��Қd�t]+,Ht���Hy�d��l��P0�}]p�܂w����cy�'�e����e�R���_�z���7Hō��` -�ֿ���)-�]����p����*mS��f?N�ڴK�4�S��t�X'b�h�����f�5����E+��$J�" �D3�!e PJJ���9�ȱ5�|�P��c�۳�&0H��� ��8�Q�������8¢S��1Р��(��M�_��Q`()�F�u5�/�hի�ڻ����=y+V�-�������4b'�_�(�%������-���KuRѓ������c8�u�,(��&�	e7R��l�`G$���������7����5���L	�W�'�<x}�^�z��N5�牾f���M>��0��W}a���4���fViCiG�F ��n���b���ן�-3�?׳
o,��g|���{1�B�F�Fh��|������&�[~d4����q*�T0?��L���i��"ddT���'�Q䞈ӊ�Yb{��`RT/L��Û>F�4w���p��J�:�\�;��dO�m����M�Q$���uţ�I�����vĕ
��Nf���̉|4��s�ڱó�Y)""TC�&��[m�،ђ��Q�j�s�E�WW�0��o��s�6=�ix$�Et�Xŗ��eޔ1p�g�CM��]� a�s3��Q�$>s�	����.t|��gb��뜙V���H���{ؠ
�=%O>�O\�Ӷ��pQ���/����b�f�1pP<�:����/���P���6�3�����~���ƳV��$�צ�r�h���+��OZ�.��̣�����sq���7��k�fPY��z�5&�x�=��� ����n��Qx����1��R�9n~��a\m�
�R2��$z���z���Ll+gJ���y�jH����W��b��`��zJpB��m,��I�Z�T/�
l՘�� �Dߝ^��
r[���~.��Kه��[��Z���ʫ�����E��Ч'A�{�Ռ%V�e�#G��2��Dܮ��d�'��U)�/
���
�³��-�2���^L��b?�`��#�����eK���]Wt
D�����FQEbRy���	E�~��Z{>���<�T}�%�}�R�,�b��=/4���L켢kv�@��)d	�	\���C�`���e;�F�J��Ũ8mWr�/A�҃�X{mk.]@zj�_�#s��)fƬF�H�����oр@��Ѣ�g�C�Q�r��̷�qmC�b[�_ĝ蛀��X8�&!�����V�j,� ����bg�(x����b�)٢惂�O%��ڜ�+&�7�� �7�l�t�H�iQ3��6�mٺP~�� )�1^�v4�<3Ymg�2���z�w��Tr��r�{x_�����͎ao�*Is����d$�J�kD���6Sj�:�2�i�Q�z��ƛCޙw<�����b؏��@�V� �T!�m1hb���>*r��h���A��P"*�k���4���ˋ��� ���;����@L�{e��̼�Xn/�4�I�^e�����v��zk��Z��� s$;��2G��u�l�6�F1��.:R���?�hu�����c��{$��E����#��t��� v�V�ʹ�S��VIOu �
�&�t"�ё@����]��[`�%�:���D*�-�Ƌ_�y���4���+���7U	�'BR9~9�y���Ok#D�@T�fz���p_���k��ܵ� C-[�<mp<@R�$�K�Vjq@|.SX��X��[ɍu=��SG�1���*��G��`��k��k:�4o[�M|�(�Z�yj��IgT3��!�Q&^Q���ؙ��_a���L�@K�r<O���o���e]Z��W��B��o�(�;
Z����U9*�|y����2��©�n��
l"�#fe~��줈�f�߿�ZW�9�}+��u�f�u�NJ;�>�q��ŕ�L�I��3����ʰ�c�p�v7� i�mNs�da,���S�2h�7�� �� =Y�R��
�(�C������Z�O�v Ü[�ub����
�U;���jP8�(���C�D�&�M.U��t��*�aٽޟ�6}�#`���&��3SФY���3A7��ҝ���ǐVU;��o%v�z��mV&B�?�@��"b�C��@P��g�4�fO��GOQn��G�>���cT0VrR�\ُ��H����{�?BU�
op"콻�ݔ�����*�� Z5����?���1�"^b�g������ܴ�-{Ʃ!���������n@�0g�䭘�LtXi�6zǞ��[���ؖ"CV�S;�p�r�mj
<�HE�-�����l}{%�j�gz;(�f�,��8kp��U��Q�&��q�_�&둍��+L	�����T	�C�eK�U)q���l������������̅- ��*��H��Z��$�1�6mY��Z�w�Ռ<�=A��"�~�Δ�YI(�Ϣ�[_�[B�d5e��Y���ګ.����x�$����k�������,��9Zz����z[�R�l\��_�{|�AK�(R�BX�7M����d\�&��b��Ϡ{Ձq�����O O9�w�dz�
��%���m��5��0���M���(qM��&��"�|��-ri�i8�z6Aa̗ʓvJ��ln�:@N�^clb�!>sۊ�m�{Ij �� ��M
�$���\)�p���؄��|��o �"b-tk�`㗬�T���V��~�-�@�k�������Y�Gz�ҜÁ���k����(�@�:��*`C�-�i��9Ah�#��+�P�z���b�gc�Zݨ�'����"iڬ�t���$�zPN��a��5}�8λ<Aj���������ԯ��.���{vtQg�`ޖ�R���E~5���I�-��QU���0��6p`��"��&���]�{���3b�!�K��;��Le�Ʋ� @�T���'I@��%:�X�7%��yJ
|�����*�$祙�c��U<��w>�y�x�G|�N����/k@�2��Ɛ9A���5�ٱ����;��lF��&�=���R�&X�JfV���}�&r/��o�v�F!}ֽRi��cy��E����ېOޥ������u�~](z��H���7aJ��R'U�c1l�������3u���T���*�|���p�^q1\�20�P�P�4�58#b��04Uý�8M׿m��������*�]��37�Ё�����zlP��BY�i�C��K�j�z���9���/���������]�U������E��Ԡ*��?��g(��M�s�b�)��'�Ɋ7�PJb��
>D�XDK��MP���Wžt��.��'�ϒ��c_�ӑ9�N(D�֟J�sX�F�NC��'��K�-'�N��vc��%#!���Sq��g3lG�����~݄��IJ5;�Sgt�i7B���e{&�/�.Q~���@U�sl�=�ܕSG��~�f��Y��K�shw�xl���u0}�LMIQ/���� �hd~K���!Y�l�|'7��SON	NjSۣ���⺖�j���.�4|��	���g�(Q�E*~q����Ď���r\���u=����%rS���4~���� :_��Fl��X&���QĶ���Ի�벒H�	�U������f`Կ2j��:�m[�h�y�2n,K�b;�8�簢�ZS�Ŭ����]�p]�`��v�&�B����D���������P9�:[m[E�$�grnVm_H3�}H�q��A�r�hw�xȸU;h��SgQ�����͂�+���t�}8�N����A ���Ι�pLja�����c۔��i��zK�ٜR(����y��K�N��z��7���~���W��3)���t#c���-/o�Y�!��R��|ͱ/3��%�)`ػ�/��y�u��_(ą����C�2���I�{�]_CJ��PFAV��|�n2���O�H�Z�XC�i�'mh`��X����Gc:�K�0�Yh�(�f�f�g �;Ov"�t�>U�@�7b�a^u�b'��Yd���2��ig1��T ��\Ε�<IN��ڬ����6�b#+�;T$~�xB�>u�P,�#����t�nOe�2A@	�����$g��2 ����HRBh1�vF<jtg��7��F��S�0(�Au㤳�7&�!��&�X.L D����c���v�P\\�x�mP̚��^���P��B��@���_f8>�hIf�V٠Ӻ;�0R��-#�V��}�lIp��^I�,H���ߢLT��/��q#9�����s�_���7T�K'�m�1�[��������<�|��f�ti�+�'(XJN��4i	��>;�ǆs}Y0���&[Pw��:��:�or�`�n���m·t�G�6�WԱ�s�.d�i R�a��^�I�j�Ư����Z�N���qe-�7�S11��\�Hv� 3���Kp��lUi�M@~��Pԁ�c�l	�/>e�=��6eSf����K䧬 �4*�[�|s���_"仝_9UK��euo��7;�����?�у���g�>�8�t�Z´��	Z�D)R�w��;'����5��,�[q�B\/5v	�:�m������'aD�]�C@oq�����(�'a��c�'�&��rn�X7�!���ȠcvLN�����֛;�sW9�\��TAL<j�1��<�t>��g�5F��� �ė�֒*sj�a��㍙�������J��	�����τ<����8����_�tk�������3��h[i=Ҭ�'�d�+�o4��o똀���	+��ޜb�����*'�� �C��w�5�e�S��| ��_���u�Փ_��N��q1	�cu*:�嘖L��5�pR�$NIB��^ �˞��(6EDĆ��	�+^�Óx:cK��D��j���qRY����/�eT֡B��X7ϗ�����t�K/�}$��e�(�6m�d�W��~\�6yHG�QJ�"�@�DK܎2H}s���n��;-B�m:Hi刑y��<��u�)�i��7����#��W���%G+��3�����d	�WlQNϪ� Ct
�~��#��[G�ҝg���l|�:��eL�d.����^0�;�ʦ�{��y�I�^h��}�$�͘�r.v�J]�B-�_��Z�Q�h�t��֥خW�ZZ#�ud%��q��фlBU#�2{�8boPG$�'����xp���.�3ţK&=�w�c� @���\w�&�*����'3�Qj�t��a���~�=θ?��Jl�t���WV>Hw+��^�<.\"��9{�F�',�d�$��O3b@���������d���P������xS�U.���`,$h��9�e��)�~v-�4G��
sI��gkm5>��~� ������u6�C�N�$�(� ��1Ǽ{+�\��٪H�-�Vp&�l�s,w��A�Uҷ(�}B��W�КZ2gx)P�~*�@�]��A�d�\��Wz3T�z�$>�nO��z#�����x)Y���u͓yޟu7����*L)���t��ut�W�KT�S1,2��.���Ly��`�6�mk2�+-[`�g=�R�yM���v��A,8��������Ƥ�\3$�u��n��h&j\��3@
n�������[���5`��, ���qq'�m�� �����b�JY�K�7]Er�+9�Ϻ玗x��n�\%;Pv�o_ݐ
��_&�^�f����hCS�*��H�C
�P�%	m����$VI��Q�|�����0�;r
��7hc���f"ǱY��u`�;�&���y�����?�.��ue�3�U\X�(B"��f��
a��0Jh�$w���_�B�W/b���L��C�?���p�U�1�|Q�P54h�5֞먤ѓ�0�ѕ�� |��������r*�Ná��U��¨�A�Io�h�چ�gMwKy�k��;�����7�YT!dn �T$�_��v-��s�K�̣�K j��窣$ZV�ܲ��DP)B�Tw����6;W� 44Id�t�~̬	�� �ors���r�Ġ3�[�:�6�4�]���[RW�hE�7�rsŬx�R����ΘDʜc��w76'�������q�R�S}A����	�*�ғI�qf}(���]��*�������t(y��Di��}��U�z�ʕV�<��L������������:��mD�9�ň������b\�r�Ș˽��cW~��'#�\�Lِ�msm���V���|�F�)�hE�񬉄k7���n�+��U{�mM���I6Y� К՞����l��r�ش��ӌnC�=���I�8S:}բ͓�Ib�;h'_sZ��sA�{r#�3Ƚ����Z+f�#�����8��Ev��@4�G_O�BŘh����~��
�<�쓢foY�����"�ѥ@���>�F�n�D.��@.���%���ɦQ����{)�̽4xH�:?}Ms����^S�
V{d�x74����R��t#H#�>��޽���q�(~���w���E�g�Z�y�\�����[�����e��N��LQ���l� ��I����1̛]�����T�~^�ཅ�f�	�c���G�|�I�D�.'Q#/���$�4�z��y��<ғLO���{��ׅ��zT�e�r�J�k6��q3�����;����u��0���ȱ�؝,��l��p	��66v����=e5�J'�9c 5�|��8u����|���kGXp�J8�А��)�
�[��:�0pn���XE>#ZWw:xv�̊.Y��E��ڎ��f9�
������c1uW�=�P�G�
��7����X T}���ܮ~������ˆ��sm�G����2d�,Z��jH��#��r�\+��G���4ze?	��8�`��m45�'2̭%`}��3��-MJ$�O�$8��?`�a8�rJ9xفM�e�K�
Hwqr�6I	�VyHH ��I�5l.pm;�15p��p��C6�2��y�߿�y�n$ �l:vl�a�m]�+�?�v�r���6?�,T���<_�����.w�۴-���4��SI�����F��W�N���S]/�h&W�%x?��zʼ�6Ps�	6���J�i=�0�}j|T�n�]�`��U�$&��p��B�o��ҹ���K=��=z)�M�+��тV*�i����!�~#���l�HaK��{�pI胦����t��nݩCj�r �X��&�t��?[u��2F����*��jD��g���S�Z|���wefS�՞e��W�6��o^��3M����
8:��D�]��+b�R�J�ڋu<���Jjñ%�8��B4`߾�)�FV�֥�A0$�J.�8:���?)h�8������K]kLRmuc�֯��8��)������0�Op�E��]B�f�Q��k�q�?
.Md��h�0�׎���7�=��^�r�aa������Ĕ��^�w41�(3�k�N�3�o��y��P��~�~��#�&�p��c|�ı#L�T`�5������&1�CӁz�h�L�v(T��Н��y@��ɦD�?�����j���?� qQ�+�ނg�}-�'������4���JcϥӲ"�����h�E��]��FF��j��L��
b ̽9���-������ʛ�����6$(�~mǙ���g�������F�uX.L�T�R��@��ai��A�[/)���Zأ�>MN�5.����T�9@�"�:D3�~�0�,�z�r˧`���H�=��2����!�ib��xܪ�u��K��Q	o*�9A|�F�"���[8���.As.ʙoxM�=�D�ܜA�#��³c��Gz�#Wi��zI��D^Y2aF`��+[�o��	S�$s���ǽ=��[��<��ѯ	b��=��9��rq�ǟF��K��j�,BC�M1�K|�����*}��{���O�\ʂ��t�E�uS:Dm\ah�Jȡ[���f����2��A��4�g�Y�������6��x�`�I��H�'���dX�}�ְ���&�`�Ҏ:E��HϜJ=��&}!hL�M�Q�y��qE�nj�����T3�
��$�9�>�ߦ>"�tp����(�������{��#ڙ�~`k��P�cj�F�x`nP*�^��Z_�sl֧	{�r�/��gPC.�����8�tb���X��N�𯵽E�t!iH��yA��D�_y?ӆ�J�Q
���*�����[~���D�F��5Nj�nL=�ȻU��e�WT����k\Y���E2: ��?��lp��f߮�����;aw"�Y���̰#���,p�rJ]�;���z0�W�|@�z �7�X�I�\�L��C��
��[Ǭ*�Nz��>�;�hc��
��׍�O_�q���٣3إ�3�$�j�;g�u$�
t��&�>xG �}��G�`�����k=���+��ؐ����ؤ:w�YΠ���"��.��2m��'V�/���;�E-�9�/��
�{���&�1
�S
E����V|%����؆e�"��>���̼~���f] ���%NiFI'�?�V^��M����ϖ�**V~bG���_�ٹ�3���#��q�x�:ӣZ¯��-~�U���&X㷏J&~��JD���v�3?����a�����x�~��r�V�������F[�:P3�{�x�q||{�`85�T�*+Fy@[9B:)��Ǟ�{����7��ڨ�"9heN�r3ȵ?��6�P�xQ#?���ܠ����B�Kc�\@"��7/ŀ�]w�f�CK�B��QR��%����hn(u��!?~�>&�`�eIJuc�M��%�yQ���Kab��X\. �)L���ݱ;q�l�����a[�%yZ6�|� J���}��0��p���g��n*�&�.��-��W����e�۔Er��.΁|U�B
�L2�z#�V��:9.I�oj��)͠K�1Z�w�tJ`B��5��O���^�Җ3��h������*���q'�!�k��eҀ�$:��Ix���'��P��Uz>��U�?�-qO����CX��
:ذ�аD�|�P�#}�FJX��HQ�4�b~��b��r�S�^��'�bX]ܤe\���_��L"�����K=�)��jy��;>IF����|��e����bX��tī�2�0���P�X�H�F����e�=��������k`��Ǯn��ل��y9��);�lB�!s�yMp^$̚gϵ�7v�5���20RY��R��l���S�..�MBȲ��m7MQW�d.��U�m$r𓤬{I`l�U_�q�r�o� ��ls��Q,-�Qlcq$���viJv"�t��%�8nLO@,I�ob.f@a<��J��*H`���.S���JQ���Ng���L�8�v[�d,������K;�T갫�el��.�	�iF���"���ęl�D��9
eڱ&W��,M�e��eh���`����x1� uY4GH�2����m�y��L��.�pƍx�d�3ۄ��n��������ż�1O�`��^<}-�C��%���s���p��3�݌�߆�-���������1LA���b2�Ŀ�C�=^c��0����AJ"]��|�K�2w�.�-����|�P��k�X�y8� �P�Z|F��8��s5����ÿ�'���=���te�A((���1���'I�<Y����I�k�nE��C���x�~G�����@.��4`@����ޮ�1F�B���?���t��Ǽt������ݺ	dG�޵\ԛ[Y�-���k����~i�:*xLC�|��IkG���@}v������'�X_�i��|��� �W�c(B}���y�XRc���l��(���� j�T��9na������ʁn�q�7	l���e�M�����eB��)7,��Ks�
9�d4K�@��&��0��'����wa�ɬ�#��� ��8o�iW9�"5E�ů�0�<�ޤ��!Ƥٰ�gK�}��d���@߀-�!�쌞H�fSe&��y���;}ѥ�@�s��i�u�L-�QOpj��Ll �Vh[�А����#"�����J�c�Y�&������b��`�e���J�F.��\��+�q�s���:+[��ޘAX���޲���Ɯr̤��n�\STG�<�ؚ��Se�\��J�`!��{��B�T�	{X0�]�V8�֤���2����k>�E�L�.��:��4�j�rڃ�ՌlLǭR�&�W��y!���ئʨ'tk*̝�td�n&����m��e���s�W�A�X����G}��<�r\���$3��}��
���Q�g`4��wM�+u��7�5sE4 �CS�_��gv�r
�=�R!gH4ev����yx�=��{gv;�Nw,�>��3#5�t�f�����������7�Ï���B���9y��3�F�`^�zT����r3c�9Z����X68EfLIW�y���A5ӽ��]��*;��̟#y�G�0=9|4�`�!vBp�y֣?��ŝ:!,���7L�M�7'�:���:�Ë�
��KUhz`'��)�[K:����Z��c<���l��ֺ<�'ǉ�9���,ʔ������MS��׎�EA���VՁ��C����FyHa��ف��ٲΪP�iP�����|��y�S-�g�{��(�n����.��0,*����a�!�ڃ�d���P¢q�?/��}���>�v�{�@�ЈמW���!dFźJ)=�q���p�l�f���
���p{�1�|��}����:�R�����SҾ�h�%J��A�����I�7P�LBa���.�8^��M�0�X�s!'��T���"��	bP%��ټ=�G��w�L�W���
鐑VpR�d���~
[�Xv(�VW,��ɓ�h�^�Ȋbz`S!�j}/F<�C���RD�4$,qz;/��Q*bM6��3�2�u���V�.��ޑmMUE���R���U[��;�́��d��NzFj%��H���ω��G����3;�;zY��vx���yxO�5��ګo.�Sx�O��9���*�k�ްՠ�ڷ=:������.��;�v����ޏ	��=�f��U���5���%���W�%��+x�p̅�8[��(X���x0���rT�v#NM�~���C�$~�3�.����B˵��8e�1�aϦg�~Ud��pE����jXA��m%�&�~�Zt�{��+�Hݞn`�f���W�/�:���k�������`c���Ո�NJ��.h˅����}���q�a]�c�,�RV���F��jbm���7k*��-��`�y~ 7�����{��V���P��Lmy
B�,+kz�<����;���l�ͯ<��,h��/m�||��]n��3�`��K���0�a�Sk�~'B,mC���`~ßBؐ7��Au���8��	��3f�{����ҟ��΃�)!�PD%oY���lJ�	*%����B�uk|�|��O�'�����i�޻ǒ��'+��,��f��m(:���P�� ��ذ��c��*�
N�h&�V�W@ d^��R��+�*Wj��o�[m#N�T��F���{���܁~��:^AtK%�5p��}���$�@;�K5.�崇�֟L{�*�@�]�Pd������Tk@��y'�?��h^<�*��d�Yú4���^	Q��PŴUEwDؤK�n�}PW�>&ۿM���H��q��igdqޱ?*ekD��B��1��8]Xj<�g0+���c�R�Yx�������L�g�"jg�c�yD�;�|�c]�ʻ�`YZj?l9��Gy�Q�(��|!���h��z�tN2Ư0d��\����������&�1�����C��"�)�]p���pg����YR�R�-������5l�o.;;�ם"?�z�
z��v ��{�6>��S�:v�;��l��aqܤǙ�𲮸��S�	�+�F��	�[T���ҿ�;$)%��� ODpmLPKT�����Qu��R�Cԏ��=i�$ǉ4��~�.?eoh�֛�1��վ>ȁ��wb��ri]Buξ� wsV�{;B�˫����
�$/���= ���Z͂�PQ�{��t'V�>*�s������LT��o��$��3V�Ux���r%m��q6C�Y�Z���O�K�*��
翸���B���Drx#t��xL[x�����\+�g`Y��uv�4� K�8�ԩ�UP$�� /5;�ѝ>Ӆn���ϥ����O�^��C�6�������g}�� �Go�K�K��L�-7c��+�J%��u$��b��3�A�cd�kɶ�$8T�28�O��ԑ�h$�a~hj�]9/Hegj
焽�:�a�։R����53�j�� �wl ���Q-���~���q��GO�)*� :Q���-&]�ݎ�;���-B�Ԇ������m��OO��N��V�[oD�x%�_��JD�>�v��v���IVR��(��o��+6d�����K�.#B?r0�����l�ag��n9��2ş�}X���(	~{�0n�p ;5���p�!*.�wƲ=t���-w�N�	+�LfNO��<m"���=+��M2������т��j��k;��N��/l,n��@�X���Ꚕ�x�~�?���Y����TQҎ����܉k��ls�t�%(@�+�\] ���Ý�"������<�q.wJ]��
:�&�i�Ɔ<w(dQ��X�dw�aH*���6�k�T
1T���%��x���jTP��x��3�j,8��������a�E@o�.�X�/{ս�,�ΖB.T\:��i�������{�E�u�Iͦ#&ݜП�G�F/!5S���Y��*�a��J���V����2K=A�fΦq#?x�mo�3u^<��k���i �%�-���e��N�η����
�m���h��z���l�SK�dM\6	r����/�]{��0�!��Q�h��sɛ(fG���u�B����+8�V�zY�Zfw2�M�m�B	�h��cmʁ�4L��8ep�I�U��|�79_��M���=P�'��j秏t�;I[%p����ꩡ3��Q�y���j��5���=~�!ƌP��XiNr\��$�;��V�B���h�7�/0�)Xq9��Ạ_6&p.QA���Ӵ-#k ���зGI[�c�K�^��#��t�:�-UP{x�R�L��C����^��C�Tx������?j}�t
�LY�w��p�*�����R���wĩ	�hx�7r��3�����]�/<0����2��:R+�==h&����u���c�-kP�8�[�)�g\����TnM�Kp��L��@�N��|�c�<k�;�� ���
ęϢ�i���I��b�OA_�.�8��� I��T>��Vd��7\'T���z��f��{߰w�¸Jg�T���7,�=����
Ip@�|��v
D�=�%����5`�b�j�8�Z��CQ�M�BĎf-�W�g�i���Z�n���� ��������N�P8�kJ�f��^����bc�]?&<_ݲq��n֤�dm����Kp�s�Mb 붆�����-�I�vܰ���xp�[[Jc�:+��)���>v���w �.*���$��m?�!ѸRC� Rp��k)ͭ	�U�f� � �������Py�2��SE�̛T$����t�S��
�e���a:��S�n(3*�!d�
��󩥛@I�h}CTA��˨�����A+��֊�3��@��oZ�K	�.�%�� �u��T~��M��w'Xx�A���$��)�@��"�X��H��shy��t�b����ůDx��{�ց�6Acm��򗪯h��(�Q�n68k�D��ô@B�#�Zx������~u�<��_��3�L!�ˤz�o~�yS��p�þ���L�!F���eZ"��fM��� ��D�*~t�bHP�vHX�|���� Ku�{]ٳ_�����H/�V�=~�
h��}����JwH����4��Q�(i�����b�R������"��3��S�}��{�-k��IS���haE���/}�h�Ҧaoq��1�1-�Z{<�A�o���J���}&��1����5Zj6"�s�ez"�#s�˲E`_I}�MUZ��wPe�R�c�8ٚ'Pݤ�V7b��N\֦+�g����`�a��I�I{tA�A/+S%��l_8mN�]�&�)��x��/0s��x������Þ��)DYNI���z�X��2�~A@�iK�-��p�}_�H�#��y&�I|q���'^���W��f:t��z}[�|��W�k�z����o���J��#K_q7a}Uj�
|�}�m6�P������
N�{�V��d�忆� �.�=�L����t�'�w7ժ*7���@OC���ϸU��
6?0Gp1�#��+�L�=t� 4�!\�[O=�}4)�`AB{�{��r��O�`q~#/s4\8֥J)��*��&��`|oG=R�#�$�ű��C�$}�r�}����.2 KPZK��Ȯ<��t��0�x�y�0�f���!8�~��Gy�ۖ'?k����V�y��M8Ʈ�][�-������D�ϤN����d,7���Ǖ���S��iu�<���0x�4س���¢��'m0�� ,�֏n��e�t>�]ǡ�4�L�9N��]I�����ĸ��Kc��Y��U`=���!/���4���� ����L!����^�n��a#��������������]�A*F�H�@��f)|�Q�{�? V�m�W���t�,q���]�< �e��^����u��2�������J�v���I�Z�n��F��� �W)�8���ؖ���`��SrJ�� eH�����	d����ǩǷ�u@�ͻ�71'I����������LJ��^��&�C<ւ�|����Xך��63|m*Uq����3 �����Q��b�Q��F1�̸:����^�mw��� qz"*����4o���2�t�P:o����>��Efp��BN����"��	�;]|�8���5j���!F���/*�(7roy�F�߆@d����=�Q��u�*qU�.��7!��uɱG�i��rL�hhO�rj���;�r!֠���Z|_��ü�A6g�yk�rg� y4���,Х�e`�C�ܧy�5Q�G�1���o(�3����*z��d�\t+����="��~#��]1�PK���	I���}8�B�CD��f�U*j����_�0@ �됆��R����{bg�����"�)��I.�]��vP���3a�N{���tS���3㸀Y�"[�J��ֵ˪'A�쥋2+�aMU�uaQ��v����mu�p!J:�AOs�ﮭ�ف�	~��E�1� lk鼝a��
�O������a}1I�L>�ǇO�GCl�[�!��5��-��3�H�N�G�Ī�6_��WA*�z\�"KR}�av���B�+}���-�\������Y$^�WK��l�}%!1ޯ�p�ÎEg$�z��bi���X�m���!X��/��JE73������Sx�I�nJ^O��p���5"(d+�i��`^!�`>��]}�Q���,C�3�%�Q�h���ZBj���<U=��|�2��X�:���h$�!u�M�����I�R�[�揆L��e��Y:c��_tD�������E� իQ�k��
�L�n���I�,�~l?�'�S������32�7B�=:X����?��!u-5TP�p(P��4&8$c+D�
^l�HG����������X
apI%LO���A��H�M��5a�����^SU�^N�p/JڵWt���ʮ�8��y'��l��+U���Nw��vX��sS��nf�{neA�� N��G5��;��We:υK7��9�X+&n�lߦ�ol��� Ⱦv�\Y2Q�*����l��C��0��֧`ޫP<�`�(;�f��}byv�;��'@?we�]��@�r��~ Mn�b�`�V$��`�N��-s�
�od��y)Nj�ZҠʫ�˂��}���~�q��g��g��4r}��s�c���Z�W���J�T�j~�P<�H���rjad�jlE��aU\���abp��5>��1�5��d4�/q�@�Ȃn\I��%0<�<������)�;���5���4P�=m~q��@u-	
//P*kS�o�&!�b��'\يY{�� ����"�8��R�K�2����:O����t��sxj�75���' �K��g0ۉI�c�SU�}�S�2?L��R/7�׫��1�F�4�4�������g^:k	x�����4�R��bH�\~�2a#$�wV�� *b1�d(����P|�rxv��T�bar����%R�J(Vn�̒�&/�`�2pܹ8��p�p�ק0�L�����ET_7t����o�Am�Z�r�O�7�Cg��e�Y�b:�Eɏ_��Lԫyj�����kfb;�2�CѼ)�?�0-�s��T`%crDYB�Sxﭜu�ª��4�����(�(�߲��SZ#I�E9���W l-o��qM,���@�f{��"�~4����_��gw�uNs�J8��5��k�vR��
�<[N�m�J�f�*��p丈���[�T���A�RJG�wӢ^S��/��Ṹm|^��V��1.��(#B�S ���B�XP.׿�B !ѵ0����±~�p��vk_y��&�\�ܣ~>Y��"LQk��^���D�o�d`�Q-t�m�fW9GI�?��6�c�0<&y�#������ׄ]�Z�����<OX�,}���is�9�-(aq�8�E"��ʋ}N/@x�.�/"����]!p�Ü
�d[�њZ�����}���ՙØX��Ѵ5��'<�v�ڥ��v��̐Y�N�U<��'1�0J��ؐ~��Vu��F�<��k_��I��!yL
��x׳���<��B����~ؐnW��B[�/�WW��k�n�.Y��/�I�jmv��r&�
I�f�+n�����]⡰����>��fHN���n2���ݯK�)��@OGF�ⳛ̨M��k��t���U�r��{�#H������zi`y�,ތkSI'�V ��w�ͺ$�(������S-T}7���G����yQ&����NY�[���E��SX�G��P��^��gg�G���G�L��[e�]}kIeb�ɒ^u�a���:�Б��#
��t�
X,(�<�@h'V�_�D���'6�!6�B�
[�T�h������wpǏ��|+��m�4���?ܡC2J:ؤ�B��;kֹph�Ԭ���)8īp����Oy���]�c� iA��P}d������1c���|��aK�(y�*4`�\��H4��>�*���p�J�
vG5�w尥@V�U�����rx�y1詄#��p^��}���L�t�ss$ ,n~��*A��5 ��AID���'�R8�i��:	Y|p��Y�dn}"�U����s��7�c��d�U����,_�������M����\�kp �H������������v(0�Mfb�6=vxZ��p�*|bz���:C�s�͉��� X���y%y&��R"�9V�����>�� �mC�:��@��a�<U6��C9C-$7W�g�Ea�a�Ov!��7U���i�g: ~"�T��3+_n9���m/}'K^��2�7>b@l~����Ю2m���b2o�9d
��1km{�, R �=6<��= ka`��~
�:�E��^`ߊ ��d�F����6AZ�)�����R�J��[��ݲ=/�!��IdKp����w���z2��n�A"{�ɨ�틶�R_��y�	���_$_�kMq��6��� ���~Y�@ ڭ�J�"���c��=�Ho��3�T��Q��=�w���uk��I7Zg�z���9"4��g:�T�԰���
����$�ȿ��ѱ�=h��~8���(�pz2;��`8P��=�qُ���n�[�&�?�әEEx׵�i
yZ`���-�v�39�b�����,է��Ka���j��;�("7���h�b"=7`D: xd��ͻ�=��6w����JSZS�)f���.9�ǈ����1x��4����5c3G*��P���jg������d�ݪ��߽b�\����'r��\+7��eȟBސθ���i�~:�r���գ����6ۻcu	UJ�/D�P�4�Kʺqz�.�Ѵ�-T�T��� 9W����;J�-�c5�y��9F�T%�J���"��l[���R�����4�����n,�=���o�Ěm�ȇ�':}�#ԭ"� �n� ����(��t�*�ʷ���[&B�� U�4u�'M���+ƀY)U�j�OQ-EH���JjDa~ #�A��X��D�nF������ L[��y����ڎ�
�LUk�u�����V%��C+����|��#�U�����>���4q�k�7wYh�@"�N�@c{��4R����cʠ��s�K�~T�x-.k����ُ�H�(?B?e�A�=eJp�Sy;&�\֐�A�1��b�e��f�ҭy�� ·?LU���Ҹ ���4�!'ʿ�{Y�e�x��~�MWH��%F̫߿8�.T���Ю���یv�G�[y��
f�k���Ж��Q-֞��˺���¤j���ǜPjS�C���e���fgd�̄ݗt��~v?��Z�v���-��p�{�;�n#� Vz5F����Oݴَ�0���R�AUC�>s���:���O�18���,������3���/Y���8��Յ���ڲ=��eJ4�w�f�7�����UUXѠs��Rƭ��-"���Osy�<��Sk�
���k?�!U�_~�z�yC+d_
�@�'4����/
�����:��[��o��W�M^δ�R���Y���4�liR���|�yx���D��J>��w6_zّ%�h�q��N����Q�ףּ�9�I*,�%�>�aW���L?���*m�,�qg���] ���O�\���	��B �MVP�v�`Ό��]P������C0��^_���r�l�1�w&U����j�?]���ك��_�$\�9��5G:�_'����ONVF6�\m�쎩>�9�Eg��!M&ț����;� ���tϻE���|���5�R����
"��K�v��op�og�N���Iq����aS	��<��P~!��PB�=�l�	�mx��@�H;#	%�9<e2㹛C�g�{�_� ZA���`�ؘ�T*�헄H�9i-�0ߓ8�m�-i���X<�]���O���haDG��ǹ�[q��2�W�}hqua
�1�A�x6�-���<jem^�*a�A���gۛ<�!�Z?Ėz��=+���2}я&�~>��]�%��d
{�mT�`^�F�G��]�)Wک��Mn�)�����%�e���ю�ږ���$`�'Y���ǝ��
;�P�� �"8v0�<��pP;��d�cClJ~��qSQ��:�\d2]��j>1�H�ZO>\z�Ck[��� 5 ��<�J�^^�:h7�	5?�7~m�,���*{�F#�Xf���L
[�ZH����o��!��I����x�荻���#'�
K0٩�_A<�(h��`�ԫ2߉�<<�)�k	�b��$
������T%f��3�u�5�44V�	�Y���x>v�q����W�R�[���v�1�T"X-"5n�=IK>�M�59�V�$ul G�ٙ1-(���,��mSUׂG8M��5)�aU�ϐ��	'3�w�՟�J��H��gE��^���А�g�Ϥ*���6~�0
_͘_--ڐ9�n��%W��&D��I |���p��E߲����W�z��)�.�q���d���thh=�W���:M|�j�Ry	(���#�Z��v7!�}���Q����K�?s��>���F���<�Uq�}Z�㎶u֗�	w�
�1cir�x�<���R7�C��8m�_���0LK�0��8H��{�p�t{�*��\�Z@�U����+u���W\�w�����R�!f;_-T$,��k�����%߰?�kI���߬��|�+�d�m��'2���c&*??��|n!�+I�n��z�B��g��p�:�h�`A,�+%��ĄZ�՛o��@�6�kS�Qj:;ΎMԒDKZ"�}�:�ڑ=��wɊ��/�5��@�"BV3��nK��1��B4��$:��yf��k's ������k�W�R/�l����0�뽶�+S�����F�R��p&v�ͻ�T�`}'-�O�⋣�4N����"x�Xt���g��~�o�\��`xZZ�,��b��C��e���~��ȝa�M�:iQ��F=���gu�T�m^h����x�e����ݒc4M�)�j���K��ܗ��Y|yx�f���=�F.t.�J�v��r̡��E����˼�O�H=ek��E^���Kx+1��Kǃ魽a�j��<f��x�V�nO�{ ͂���`�O��+���|<�v�M����^�0��PKf$i?��R��Q
΂�S4L-�f�{u�23�[Z%�Ւ����mAS)�dUOe�H�"� �gA `~-�.�j�
�HC6Y�+��Je�`���Z��B[��=WP/�L��{Uy�*������9��.-���f� �.�n��l��î-m�Á	2��9��]�+�9�?`����]��I�`� fg��e��.�ʁ ��[Ϳˆse7��w�Ώu�#R� ���lM���x5�1�$#�)`��|��K�]����kDI�qx��������9u	���k�N�(�Ad���z�������$B�S@��N$߀F����������P{5�$ u�Ϥ�H�9����M2��Ȝ5�q�^�-J0ۢ$�$Eb6��3��B�}��g���~:�����]M�uc���&��:�Iƛ�a����M�A?wƨ����k�J��R,>�p�<Y��iBQ�A�"�ʘ3��J"�&W�hP6�/�n+�ۍ�6�]l��/۰O��[�u
QI�O)��<��d����vC#(�5�m�ٸQ��f��-�Ca���h����>jЂ��X.��������;��=Ӥ�J�7UɊ����s�K|Ղ���t�0nרI�J��|�e�����VsR�Av3�ٚ�hͪ� ��(to���y\�8��$.2Y�~��)��s�>66jQrķ�M� S=�d��;w4����l��q������q��>�FR��u(Ĉ�C�}r�2���VZO��`q��F�_�4����^�j�}����-̳3I`�\l	�Ve �2I�":�\�Y��7�Xy����}/�a���#�JB�<�\�y��%��7�L{��AB&��G����Fg�gk7�G}�b�#e�J�E��T��g�ZZ��Wks�IpH3	���4��A�.�~�Dv�AK��\��Z�kv$9{�پ&�%�oS&�9�ΪAEq��?ȕv�� J�����zZ�-�l�m����#S��� b���F����/A�&�hy�ɣ��l"��G��	<Z���%���wG�zm��/--1�V�+ҳ3l9���i��H��k^���S��@�Y�Je����~�|#��H��.���3C_b�lk�z� Q)N��kG�b>C��Ă�5����c�Ў3q����c�g"��T�]�
�MwA��J�B�?�f�d�g��2f�"��-�`��aw+R}'㘤���r���z��bl:k`�C�p�K��\�_gp��K��7�(���<���mgD���E��k���z�W�#��0���*�zB�����'7�e����bK,N���裚���8\�14/� ���`�Su���wE~ Hc�MB^��[�)!HZ	�Ð�uWQ�e������U�g� Z�|&�!D����u�غ!Tn`f���s����]4�,�=�-UoA��/tw�#�Y\�U�gN9�b��VV����u�I"X�y-�ϿS���E�%���:T~36����f��=�����Lr"�'`����W�>h` �c���Z�u"⊉�?�Ѫ����D:�N"��w�T�{��ts�шy ���D�I�:I����ME�Fz�OX�_ّ����\}�T���4��ftx��XL�:i��/I���6=C �I��u+&�k�m�����p��D���ק���K,`R�~��ty�Z6z��(��꽚���y\T>��xf�T���3��\7�9j(_�t�`��b��*J���N#��ɣד.Z;�G^������p�M$�:�ޕ=k�y�?NcZ���'����u$ؓ�q�us��#�K,����Q��ŕ t�b�m�mF7J�x�o�m+n�-��4���X��o��Z]�.�&(E�3a��FB�����H1d� ��%[�D���(��$*g�
��K��C����st8�Y%��V� ���~Z�T�����,�Ǟ��t�c| ��h2����v6���,N
%��f(�N\��F'��O��S����}t@�!��>F*�!h)��Pf28e4�������F���@�H��>�Q����M�ko���C����M�uv����?��\�[*�VF���落ǐΝ�V��	Zč�-H?���t���ׄ� �|�Cpֺ$Ls�S�۪��k��L��5�G��D�Y?Ȍ�#��=���(����j!)�Q9��v�;�^U�}8��/�%\����v�b֓���̿3X�`�ǭ��?�뾕���8��M`H�h8D#��t^��S�@�٨M4dT�uRނ�N�L�3�YȊ]w���Q3P҉r}����A�oB�������^�� V ;�f?�u_����aj��.1t��XR�uR����t�/��n��o��㉺�oi���3Nʋ���Z0T�p*�5L���W3 ,3)���eL#D,��_���P1��޴8�k��a�J�����<�O��dm#�	ҍ فox�i�*��@���޳�|��4���:�7 ��L�:�@e�N_)���J+���ԳR�<=�	�>�Vش��Z�UXb�)4�2�b�:���)׼�튏�c���k��^z�ΰ�@���W�"���]ԄA���`���4vs�@)wް\�T_P$�U��{q%���0�]��<]��9a�;*;Ў'�2��5�Q$�-SN�яWqrc�J���e/;A^,};��������쯱G���?T�|�J�n)w��~�"y{�dx� cC�����|�tYE���	3��t����2L|}�c����(�����TC;W�1��ɪ8B���O=�����i���QA��EV\�r�4-�z��}����ڹg��c�R�����&#��7����Db�:�-a����/�)�a���D>�)|o�?�u�������+m�P���̓:T&��:S@1O:��u+�gޯ��j�³����U����R\F���GI�g��;���s��F�"�P�#��z��K:�SQT��j}�����{��x���"�-�����.�J��gLx²H��Z�8�����pdN��{U�_e���HV%���u���n�fc��B�XJ�C*��^g�_��E:���=8�ўn��yQ��G���5ǌ�Ŕ�iӾ�'|R��m[|z,����/v}/���6'��PIĤq����E@�j5��#Z�[+�ް�J֭euh	��t��V��ݭ���N� ˤ����jև��QC-b^�α�\Q�ã������:�mqT�>7���?1����c��m)�E��1��5��/(c$��*ٱ��{X���H�㩶�wd��e��-�_"����Ly�{��[��|W�hϔ��4�`<s�gNf@��>=��(����
䈃~��� Ώ\Q������'=p`$��X��[�����c�E8E�;��G��`��Sgs}䙳����*]jx����gg����n$e�Og��A���s=����7'A~�LwV�x<�m0!�8���ߔ�;��`m���s��vl�!h��(=��T�P(.�G�:..���y@=4ed��4�Q��x����bu3�$NLKo�@Y�H<.qN������(ێ��7�9�����8�:/��v+'|��ܲmh�[�y�*��R��$��v��X��-О���LүyQs���)�Q�mj+0�)�`�������y������m&��|Ha�n���Mr�����;;��~o��ٻ���8�r��z�<��ݰ�Z��D���mH�S��"�Fȼ���R�f�[\�.�^l�b�Ni &�����iy�p�8�d��@���#�B]�/���#�"I�7�Oݶ˭?���H�<n��02�֟��r�ե�]l	����.��J�RX�b���)	�%�x]����Z1��7s*�CS�k/�2J�}ԇ�(�()�o,�)��b��<4@U���c8˷$$Q�u�BZ��S�_/w��x�g3��*����m���?ھ8�,�t\-��(����yX�H���*d��u�+u!�`�R��V�����6����&��01�6r`2����h��m�iB��
&�[�����A���������wґ����$�?��A)�䐪D��Y筵� f;P��kv���3��We�'�k�@�ؕ�i����$�pX?�Pړ�������S�2���Uao���8`�V���0*��?�� ��4��a����(����?ډ�
Fkh,Z[�Ѐ��F򶔋�����ƭ���n6���#���~Js �l��ħH�������=����_�t���b���l�k��q	_K��E�Z�,��OX"nȲ��N�
;b�	�D��/��]�[7H���w����	5Bbv��Rz*�F�������X�:#����2V�11v3���V��k�LXF ˗8��	F/����5]i@�wۏ��|�z��$���J׶�4Ԝ=�PD=kk�!p/�u3ob;0	����$�"�,��a�P�r��C�h*��Uq9�Ͼ���}�4ۙ/Q�Lk䘞M^5��*�����_�E6�QAc�-zT��e�n���[�?�q`��0TU(��݀��Ht:��"�v'\R�dH)=_
��D�yZ�"\��N�s`m�T��>�aLk�Z?(Z��Mˣ2�l�5]���NqQjfGw��>�,v0�jF��iH?�A�?�$*�P���gc8J�8�S76x�Y�̏|8��ku*��F�S���|��/+��yFK�:���/֞��e�O2�ϴ�3S�TF�*&ãv����ZTE���@9�[״ËW��F8*�t,CT�~�ޣ�K�⋠�	3����,�1+nr�Ѫ4f�2�w�'�H�����͑�����,Xw}l0.�A��Nm��p��"W@�wef����>Q�h��a���[?̇wnC��0$\	��@Rfih{u�l��{ �nB���x{N0���µ�N1E�S�X��a��4UCR6�u-�攃�D�jP�_����c�2�@���[���_9ӎ[+�F�-	��d���Dz�����rd��>^6�e��4;q�*`�.�탲+�lo<�B��)�w���$T#gQ��c�`m��B*
�b��H����yd;.+wL���	��C R��c�{�a��\��_��k[fr�
���rͳCg���!E�f�*'e��<w�}5�jG�����v��{�u:jQ�s�������!�?��x����u�,��n>���ko�g���ɪ!K��V����}ǘ���စn�l�Ɲj�>x���?:BōdS���v�����MY�yPJ&��U��oN"P���e��X�t�(�!zt�Soq"�֛�&�k���X�+X��ox���T�!� �H��E��՗Ky��߅�e%����M�/�<�՞�B[�j\w�ڡs�&��� �����Ep���F^����sl�~X\:�DEn.��������e5"t�e�pC�{s�a�l�OK����.��U3i�w{�L���v?f��,��cׅGI}��q������K�c����.��ɇ�k-�f��󗌩�nHH�Z4v]Z�_��Ҋ�����J:��kՒ[o�6 sK���+�O��6(���,�8���u�=�=��K���$t��}7������k�4�-.��~�/�Fٮ��"п�V�k�i͹#G?�LX�	.�}<V�QF�N��oD�U�Y0a��3x��X��
ٟ� z�P�?��讼�
Z��� =SBn���H)���xwEAf��ߣ7�����q�{{�݅C���cUmv��-h�@=�QS�3Tqw����W�� :�!Ʊ7S� �r��l��ֹ�cWC7��$z�,��ϧQv��	Y�$J-�u�#*�;e�%�Fj��b� H��Y�dFL'����Hp0�4��n���D�=(�	�۬D\!*&p��F�h#��Z����|�b�������'?�9!!��a`�<�.���a3���i�-�#�_6�Q�x���1&F�F���D��>����[��Fq����,�ހ��,���N"sҘ2i4\Ie'F{�4�=������(�m����a�$��Y������S����C���Ų�֑�+ɻ�Y�����
�s���׺�é�S���&�BPgi��`Hd���g��a�J��n-��3�䦙	6��r�d}Ê���B6H�_�;3;�t�Vq�L�b�!H����M�=g�M[G{H��'�sp��j�Z���nB#����p��ڽWn���TEfG����ޛ�*:��9��M�ŲK6������־򙸫qL0:�F]Y��W��N�t5��$^R	��h�+6�Ǩ��?g^蘉h�B� ��3٣��~}�5ҌD�$s�(�`~J,�w/�>|2.�xԮ!�|ʝY$*���[���Z��![퉋�,�K�D;2;�D�1,���@Csk�$�{j�͍���Lf�!�i����%�J���c�YF�N�F	w�t�{��-	z7���1�i�	��#Z������S������2����	�L��7��x�̗Q0�Cas���z]n���|ܛ�p��9��'�K��9y��{��i  ����5g���M��s6�����_4E��[A��閾П���|�����D�v���i�&��{K�geͣ�a-�[:U�p�`��q�79uy5T�/h���c|���D��
c⑵Em��;
8���Hg����):?��G �T�X���\a̟n��p�l[����	8x�����_3�t����b����գ�i�x��.��\C�'#?C��@���
���>�ޓ��Փo{-xcG�Ru~��(���_ti8�`���C<��%e�}ݩWWF����i͹��y
��H�!��zFz��2�G���{e1���U�!��#�{�$��XS(dgs�MT�Ͳ�ר��[���s�(�c�H]L�rkV���x�a�Fл\5�G��l�`E������u�/jm���"0s�cSO91og�ŻOna�B���1���?�x]-�쁋�s6</�H��\9N�ͫ����-��L5c�`�wv�r~n���O�D�<�I��i/Y�,}�M}��Td�Z9��ϖ�D�;��0y�܍��gd'���_�~|��7�#YX`�@�;��,6ۣ���柡S«��4��f6Md�-�5V���N2�������h�9�5��]�̀P�ZJ ���g ��VpHw簽B)�����du\HZ�K�g��s���`k]>Qm���{ԥz]������5s9��%�8��d���b�������0/���w������Ŗ�`i�4����pu��!�6_�@PsзfR6�3�yAخ�,�?�6��_�vꌡ�|�R%�H�JEŷ�) Υ�c������1�y�?r�i"�3<-0x�K'��������G>��KV\x��\����v�G���
%�3!g��.Ǜ�i�ˏ�F3,��rV�Ȏ�X*rUmUf"���.�hi����a�6C�J�����"��b�AaUV�[�luv���O4!�!*���ʍ@]��ʃ�FTsmC<����X��oR������)5\.B�@�W��o۸���L]���]�[�?��`�N8_�o�ћ,SÛc�^�����u� ۉ�wi�s��v%�%�@��/�bO�i#��l����x햻�~��0Ȏ��[�X�}w9�d�Å��Ӕ���������g�z_S�:������<���<)���Š�H��(��&��h9�<�a�E��1������	������ݡ��r�<3��ٓ|�yT�>rg}� ]e?��-jCbyQ�/���!V
�*��'��W�3���/Գd�1A�e�4МǑ~$�4\�C���WR�Qn�O�i�s�c�$�6/�vvߨ�$1 ��3$Ɉ��'z�IƜr���΃���@����4-�����{�B4��z��J�@P͚Y$����W�(;4����u� �b��[;*��?���Ư�!��SJ�l�ҝ�* ��L�7������WS��z�/uT!���@�������].���4v�|�Btx���8�+b)	����[,�$�K̢���wʯ���~p!�\`��x?L~(C��m�RS9<h��s�"gʃD��T�M*a8����#
'=Cs�t��9�}7�#�`��X�>���`�W�à�7@w���oX��7�zO�����LŗAxVRS����>^��D�@�=��T�;`_�Z��6ɘ�Q���V�>1HQ�
G3(�a� ��U����$l�S
�$'ŮU;6�������]6��è���B�p���¸�����S�mO��#`e�Rr��^�ǯx��H�\��0�l���z�N`�"�h�����,�U�$?��i�/�&{g?�i�(�,gwIC�AM��SQ�xN��Gf4Zz��y�E}�;���6��O��b���7���s�ǂSFr��1�yـ��%`IQ��]�*EDƑ�tr��{�"֕�=��7�;p�ZmRB[FY`�_Oߐ(n$=�)�YƯ�R�����9����z`�b�0��>o�y�.�w7�0��|P>��^�������i����~?W��9Y|B.�_DZ��"a�#�"'z�ߐKbu��e+N��]�p$�6�iB��S��/L#ƃUIj6�R��3Ɓ6�k��8?����m��hC�Ar������v(ۀb]�v���0�w�T�(�X���_;9V��z!@���e!�c)�������\{/y���U��`S�A��Wׄ�Z��U�7r�,Gb�OB��&���
C�p��m:�0AR��%m�B�j^���\�3���"c�����{��uX�?�B�d,�^3�Z��"[�������,���S��E���c��׳WX]�m[E���Ӵ���ԁ�ڶ����&�������������ZQG�WhUhi��gNE��Pw�}��՜`�W��-^#Γ��~>���W�wk,d�9�1��.@�!}w" p��j�F���ա�����u��6hޗI[{c��05�sv�_C"M����߷��=���~�>����(�7��Q�`?��4�OJ!��E�.ie�1�t��a��%
8�OA*����i��;�Z��J��Z��U�ߏ���x�F�N�~��{wa�=� Ie�v��S�Et�(l���Y�C����-���d��^��q�$�؈R����(�!�-]r L�������8ۥ�M��ZtNr��qV�ey����;���\����1@�bx�}���}�VU�\�8�W�W0��Ӕ�cBY�^�Rn󭰋_v����/_���I�����٧?���-C�`<j�
a%�@�q�O�b���s/������@�	�7�7_���`"���r��q�E��H�jp=ރ9�+7<�&����j(��4��!�F^�����-��Q̵3њ��*��}�q,V=����T�Y�4P	��4i���q�����ׄ�$æMnJJ*ܴ�rI3�/Y���0f���A�=*�ͬ&����[���Hm�7��������&�Ć�L�p�(FA�Eݸtd��c�[�=4R�H��X�
]2!��E��^��l��S�#xہ(���%Jn�v���O�y}LU��ժx	�1d0�j ���B�3oՑ��r�E���3�;;�Q��>g6���Ƿ�S��\�D���8M�?�n�8U��X:K~�gW0��|����Wϴ}<�pQqȔ9�<����N��I)�Ȁ$iG+�٥*���p�x�y��:��G��*�Q��d�Y���}�U�g@�kgTV
���Ym[�����e�1�&	�(S��
`�PC"xXl׬@F�1
�
�9
õ����d��gh��0�U^9�����Wv��@[<k\a�������%�>�c�GIx
��1WD�	���s��S���wEwil���3H��6�<_��"88�UFu�V%�R~	��~Ե>(����A��ݠ����P)�����eܓ�$
��&���Of����+�.|���q6	L���v.UzW=O�I9S�>%�l��t�_�e�	��n!M#qX��}�> ��6�����/1ts���$��}�� !����X#����hf���̌��o)��5\$C&P�&)!Pe��c��(k��5�Ip��w�
�����2K.�Hi���4�U��x�S>���w�Kz��>%���ƞ��,�	՗�%�̭��U�^�+e��L骱(Se�&e�p��� ?ϭ0I�զ��U6&6���@�Ө�Fm�n=�ٹ�i�OH���"����N�>z�R�1T��R���h.qup��֑lIg��jf�������3�\�ŎUB�jUd�11������De�xS�|*韡e\�F������ъ�\��ݠ�86T�d|���g�W���t�vY���G�S�r���b�V a�.H�%\n�����f�YSh��D˘?��`�X��O�)G�t�n�N�����<�z�8��h%��P����YY��_��������H�i��Z��lv�f;�[r��VT�@�!�)���do�F��)�B�|G���4������k��pӦQ�o6��5!�q���Q����aA��d�D���B���Ѷ����`����ht�����A��/�;�4F3P!耡U�yՀ/�X��K%nw6���?�*��2@��(�!�bC[�,�^5���D�(���u��(�D����֪͟�Iǜ�f�|��ė�X�{��ܜ-����GK�����/�)�U�Yu��Rw�d�}I@bEE�����`��dZ���Y����7>��ş��ƤU�r�ez�Q�^ɮn�,�9������xÒ�ƒ�t�wt��H�2
�ԍ��.���E�J^EJ�n�K��yq���m��nD�4`!��Δ�3u}lL�
���`�Q�S8�h�Q���)FB�GR���+ʎéf|N�ÅbB�j/�߀��^k�u���J�	�<��{c�j�}n���)��X���y!��v��(ߩp�g����P�XB>�����mʉ��,UQ���rz��h��둀A�i��/K9��Q*ˍv��M�.s�557a�����*��`ӟn����yP�|�ܫ�D���ަ��;�zR�6Y�֒%3^S��6ֳ�^�p*����tiaVU��⎝w)�������b?����~�_vȮC���i�&�y9�	d��<����~���$gg)����#���_ͅ�/��ߦp>��Zձ�b��33ӓ�iJ�[u�X��o<c A��;��o!L�v����c��>ԜB�4|=) 4��%I��(��ؘ���"0,����.~am�O���۰%�!��ݜ[���./�:�5q�gA1&��<��*����N�� ('�{������S|��5=�2�*�Ţ��$��R��T
>Lw�ҡ4�n���t��㸩�d\F$���r�o�,�����ÔgY���Y���8��K��-��Ga> ]���X�gMf(S�M�9�>�K���+���l���Cd�M��/�I͋�S}�g"��r��<m�ls�D����+�V��9���=�-�{����*Ÿ@V��PJWѪ�`5��u�~�b=3'c�aFף�eC����L��J�[>���ֵSg��g��=�-8�K�X�V[-,J麈��a=�����j�|\���Sդ!�KbuOo�6Ow:�9�>ܓb�6���\����.!�JG�[(��y������������5�{����q,���.X؆X-,���:U� uz�'����C�瞪2��x)
�; sȷu��G��b��{��1!!��h*i�O�B~f[^����G0]f�¥���sb=rn�~�A?�F8�"�Tz��sy[	�b��b(�$���#˳_K���e��?aЈʄ#�E��r�0KE��~́�Wy0jo7"��)��xO��r���V��U�yٜک`��7Ӷk���,jX.�x�� Pھ���`�CP}G�~����A�1��
�U�C��j�b:��2Xq=�0�:�o�듰�mF��,+Z���
'\�_6{q�%$jf!��Cv�S�UV���Ab�`��J=\��ߓ�v�R7�f�wT"O�F� ;�3Q�_�	�H�dm��"Æ�2��!����k�����#Z8�e]�/2�_�R{��LH�!��w
1�)�?�/3b���rqB�B[�F�U�o5G\?���z#S~	��/#~�����R�юЉ��rU#�^}$�'�]���=R>����Xf����LH�{R�t� uN�~Vb��`�>�*s����xI�;�������f��F��_������T�@a�;��u���s��1���-�r�F�׀��$�5	��w��2aƇi� J?��i
ȑ�._�x7�^�u�8��G��+�t���f8;��>-��O����)�Z����%#a�B/�++ԁ�Zb�G5)Ԡ�5Z�p������C!x�tj����`�ټL�� �Ϲ �S��b._�O/�SܞV�Edw�|F�O�P��C�l5�ǃxx�Ŝ�����Q9m��ǂD��oa��0�n�P�e��� ����&����/��I.�Q�#���`
X�TJ��5U���1*�D	>� E7�<+{c"��r��M��nG/�O׎�7k��ah1(F�C�h���r^6G�ۖ��!�����sp� Ȣ{�1����
	��48�4n��M�N(`�*��2)�%	=��ܢ��I�i')Qڈ�{/I2����f��eo������5�ԛ"�Y�9X��1zG�	N=R@����S;Y�2��ī5��'UN� �Lq�ӵ��D����
< Z�6��1��2�¯�n��B�〕��X���cC�����OR��R��}�x8Q2���<�k��7!Zh�������F.�	�28|�f`>S8�/�	LCnM�_M��d̐sL��+nwy.��e��	%�;GX�Э�{S�h�@�/��7��7Ó��g�d�P��}��� �쵃 Z����5��
؆|?���=G�08�e�s�B����fTş�kJm�y0E��B^�5�A�9��\j�\Q8�����š{<C��������Nh�� wN������ѭ?򋝎5����1߇0�����'����,�d2 �^��(��0a}�]k�����vk
�o�5�T��]"���a��J鶭�_ǣ���40���=�
.��.?mfhz�{��o��ѵ	M�_��3�>'ܶk�7�%Ë��Q�'��@:���ܛ�����	���.W�MG8[E�)���M AE����)�R�P�s@�_� OZ����D�4�C&��]a�CMc�
9�{�SQ�H�W?���c(c���o�J����'�!W"�n�����got궂�VG�,l])?�GK �y��;������r�L`�@�"9�L��{fb
�:��ڸO[.��r�H�f����I�ڹ�I樄_�d�R�8
�DL�ă9A9�U�@�֥��eR=�d-��-�Ʋ�6�C���v�9��(a���[6�|� �Q������e�3��#�=b��\���:�T�����!S��ɼDN�� ��g�	��0#��&�����]���ud�uJF��XM��(0�ΧV��_�:|S���W$"|̖�3Q�1�|�.�E�K�k*чxi��"���·jptB��6\cY��0n�`է2_��?^��6[��L8㌋�+�����']��}��A���b�dB�2�p����:�~ U���y	G������?���aT���r�x��6���� �\��E� �����4��9����/͊>�0�A�m�`:�rܑ�m�2�wQh�4�$�6X�p�x����\�^�W�8���x;�ȑ�?�o�+b�k���߻�h[��k�
�ᛝ���P�#�
؉%��H�]߽Q���|��[�+�$zb,z�bC��Q?[��M�����xz0��E�ƃyh��>\�[�t�2|�*��[Ύ$�m���K�P� �uQ)ԋ��S��G5Q�Q�(qN�{��¸s�?���i��"�m�-c����- �I���ϑY�T�W8�Y2���;Z�.�p1:�P]�s媱`\D�g]�`�w�[cQz@�ǲ�Jϔ�s���$�����-RD�76�f�C-|9�+�$��I-wKq+$}_V�l���\�g�Ф�o���W2��pi��I(gXt����C�O]2Ea8�����ۗ?_�\O�k!oʺ`gU�=�2��V�\Ղ�p�/��f��u�T�%�����2�����4�~�eK���	&7f������ԝ�ngP1�3t���o��H�*HH��24x�����,sX�
��,�s����F?x(`k�! X-�ziT�S�o�HE�p.��
QD�8�&gؿ���^�J�l��_������Y�3� Y9f��uY�YJ��������V�l]Q�&�d��t�U`x���?-}9�^���"�4�w>��q�l�Ea2��Tq=P��#^�l���u���:�Q�~�
�3�p�m���nyyH�?�A��g�M7�+2X��ߗ�a9�.j�m�p��V�+s����2y+�UP�A��w���>�x� �+`Ȟ���\i����-z��5$Ԍ�E�{U}�� ����Ey�4�>s?�td �[�P��A�����U[a��T>�2�/�L�|��MIj5xk04w����1Լ�*Q��.�p����\��B�9S[�����č]��������|�����k��ġ�}F�bz��EƬ0�7��ޗ
�s�r� �rMKbj�E0��~����&�o�<v��?e���+���!n��qVFG��Dk���]q��R ���J�8(:����_3|r�(�Fژ�Z�,���v?���Lp�SR%�����i�Q�>���"��qbS�������kIܻ+ö��IZ�>�����y��2��AP1��ÉC�r�{ۉ�.�O��<<�,���O[��SP#ͳ��J?Ց����~|gO���6u4-�.����+��"g�^z�9�[��V�|�k������ޅ��q��T �陥�aS#۴%�oapZB�ZT����8��;ʌ�x�J��\�Q�@�q��.Ϲi@݆���ctc�n���ZK�Q��d�QH������i�q�X�Ћ�?�"��L6�$+����Hc���� ����F2zY�2=��L��O�n�%f"m���vJ��u�X�V�T� I�:�/*\3`8-=���^fl��#n�?�3|�D���0����V�� �h2�3��r��O��
�\k��p�P�`#j�t�c��c/���j/e���� Xl�^D;E���s.o�˸$�lI+q�@X�5g�6o�?��h��( �,"�P�z<��Z��$�V^~������k����Q��+l^@���Ϛ3�
%5H� ���!���>�%��N[[_���U*�G�/E{1��*���^�L^���AϷ�θ޻N�	���ܝ��zW�_?�ks���>�$�����k��G:H���op��F�x��8F�ŷ 3_�\A4���Zo��2�}O &\��40�O�F������B,]���� ��l��%�i}�+$Vo"��S��N������c���ՁIA�9xa��3]^J)��b(C5!�+<X�tS9-�V`�B��xX�o��3��%�&Gr��W�'����:�FE ` �V͈5^۠��F۬���q�W�	a���^���X�Q��Y �'_���v��Jk���)=T����`I탽��\���O�0��H��i, ��ԏS�8$�A� >F+���P��뵞{	^��a;��
�{j���)!O��<��^xA�:ƥ����ԹAt|��9fY�U��`�U�J˘����,k*�e
F���	�F���
�!���C��/[�?w���\�le�|ηa�u�3O�Mc7 �QZ8������D�Q��4��<a8�hD�Z����c	it�k�ɡ�Ud�g���펬�p�N;�w�$�Dn���P8x>�;B��>�J�����h�/�E�L��UH�C.ځ��Ȯ��� �E��K,�TK���[����낷��5�z�q[��^�U�ￊ�c�Ȩ�*��
_�����&�	2r�3���E:��37^�=�qMp��p�햕��2`�"Eѱ̄:͌ ��a�%��h묑+��Ǜ)]%&ci��yIt���=��<�ڞ�Ș�	`W��Q�C[�����@Ϝ<7?�a g��86��/� �U�1����z��ZM-m�,N����d�f&\>��؟���6��vo��S<��:����iZc(=�"��9ԲrA%�¹�x����I���8L3gv��>�vlN����5�B �5�l�`�i�<���oFWEp��&D=�~�u�=/�	����� ׋�P6O ��M�'�$� -�ć\���<�O֮S���N�����mU�- �P;T:p�����>Q��`u=���na�gG��W�3�u�_v��1�I��J58�Ud�&E)D������s4kփ��������I�h+�*o���J�|��]���mK4o�`���;b�z�oYi��@v�ʉ/|��z=�H8�G{0��Te�3q�����0ܷ{�X�LbO"&VwÚ{kp�c߉�<G>��>xT�=(N�w[{�VÜ��������o�E?�+2���>]��.+/bzx�4��6.��ܢ@�%���:�nz��F}3��s6��|/s�[V"wd�CA7��߼�7��J:�1o:'^W�94A���b6 ؒ��С��v9�n��4�/\��#�.��%�����"�����?l�_���\�(�D
�m�nK`d #LV{uJ���S�����Q+��,����$�`�ꎶp6��Suj���CbJ~���q�����N���>�]�68��]g����of	Bl,(��.Q���Ȕܒ�#��[�7�}�'�$��FQ�lhG���8_�Ձ�V�p%= ��VXk��i��	�e�$ȅ�!�OW4��Eg�$��Z�������9�r��(T�,o)�B	9�+�<p�h��:]L�q�`P:� �{��t��+���#�<E�J���p�e�l���Gez�(N8׽�c�$�+���lndr�׽��(�&���+`~��JO�TQ�ˊ�x���7�iʀ���Id�%��:��=�~2Se�����(�|��i�ߨj�7�� ����,t݋�}�V������)�	B���W�!|f]������&�FF�+�O�R2W�GT�v9ԥ�n��ָ`��g�s�҇���g�e�d. �m���
E,�@.}D��q���@�~%w�$�5�Oi�$�I>k9	ӬO�lC"�(�P�[d�x�5��Y�+ZDZ�B{�E�	DFد+z=���~ "���$��� #�V�}�F�
�[[��l0Nip�̿i�֯Ȫ%Ŗ������Jt����,��J[$؅�x�-��]4f�����W��}_E�ѯ\�K���r;OB l����Ф-��%ܦ��k�O���m&�2�������lT�&C(z�5��d�d��_pB���yg����]1	�2y��q^4���:�}��svk0�Ν@sohܨ�ԝ�38iP���lB&(�w�����@�a��g�<#0��y'���/-�-a���b��G�8��+��(�.�";����k^'��:��Q�g��!|�%W�o���3��H���C�6�hi��f���i8]��\s���X6�40}1`�_.�^HO�j�^���!Ϟ��4Zjў����V�T�2�3��S�.h�G���$��G�a�v�I��!�3j�F(���"H��:�A���Y�ߓ�r�v�����5��k�W�a�4�gB1�JP+ �h,���1��-G��;�
�Ov}}�Ϡ�乺߫ߦHb�G����2�]G�8��[Nhʿ'?�"\a`�[<��a�Ӂ�^�+#H/H��֭x:�<n��@G,,d�����K��J ��>�Asya�Jo�D�h�9�=Tݚ�
s��=�˺q�o�� 5�!�[��x6I��쒅}�g��T)�����tA��V�͸�y�+�[EV��������xC��H��@�C�cX*}�TW�)��ӵ$�D�iK�9z�ɤ�C�$�xx�k��ln֞2+�W�4/��د|���1.�]L�(\���y�T�� �pY2�Bc��𽻠�S��F�����B��� �����]{�R"ڿ%��~ x�Ww�6�`�lmG����!#N�\�����V��v�,��w�D��rc� ō��H��Si^>�K���j50d�U���/�D���פiG�s:���)'6)�T@hG�#G�oU清҄�� ���Pѿ�g{�8%�)�O�)�x�������0�Q�ޅ_A+�#��+��U$5H�N?�,��7.���6��_���1���e0��%C^�ݏ�����ڞ�Bz,q�d����������$�i�T_�+Neu�v�A�2��鯬{��u�-[ @��m,�H�	����J'(=��4�LV���ת��(�Q�)��X�u�o_��!ZGA���l�Y;Ē�M=�Ȋ����p-����9/�
P��|	�|���?s��觌�eX�		s^�������|!�Nӕ���$�	�ORlo���-͈`�풞oʽ/��=|o�@S�S�����;�E����?�7�éj��Y"3��a��!��J�f��؁�b��hB;�AGnZ�ZJ��(���f���'!�_r��N��7���K���2��ܲ���~ŽkE�hӕ��������C���-S^�k��a<"�#���\��_�J����LHK
2�JƼ�Ic�r:�A���s
+�X�+������W U�jO��s�is6U[���&��M��
��S=�^c�8Z�~��7����.D��c�c?ƙ*���09Ҋ�ľ��)������w/Rj*C%d�i���ì�gC�dg-a Z4�	�t���¿���a��Y�u9F�Y�5e 6O��N�{��(e��	]�x���V��|�
/u�YZ�勡5h��ʃ�Iٹ�>2>s��H�諧�`��l����2�k�dô�i-E����;�(d�������/��E�k&dJN,8wJ&]�ߐ�@�'�Qpn@r�8Z�qd�"~r�#I���P��%?�m���0Ĝ�����D�������e�x#
��w�Z۱�	c�˿�>K�����)_��ΰ� y��7���}�^�k�0�>Mb�E�ߤ�}�گ�dQm��,߃5���Þl�YJP������
w����E8��$�[����AA[�����d�A���:ʦ���Ę��zH��T�y_��&�R	WN�B���/8ae~=���]
��g�H����B�(�|��4�s
�-�q�iJśȌ�R��	emP{rK
(XP��b�Ԫ���߽d�g�s� �m�4����\��?=�E��h��G��q*~�l��@�d�G���w �s)>C��1�W�ɖx������ܴeD~�w�2Rgd������� �8�]*%1k��p��n"XgJ����,���/�O� ӭ�$��0?��=h�O���d�Īf��76�����f�u_m��m�Z��#�ad������ĳAVf���#QK9^�]}~�TS�U�}�����57�у0���8�8-��O��J^@��B])�zy@�����Ȣ �wڥ���ЍR�5����w��)��feH)��r�ՖRl�H��k�xַ�Q ����z%u+@�`i�Q̕6�_$>�laZKہ.c*&���^��R��n�Tw�<i�֡�)��a��� ��3�K����$��E>��O	K��/C���`갴o�az4s���X�;��#�7�W�iB�du˰1(�k��T����^=3����;�պ�\�f�(�['H�lp���g����lL'�R�k���8�,����k��'}�W6��E�N�E�St���f.�M�����)�* �u�����p"~�r��D�w�[9ՔreX�Ɏ��sdf�X�e���I~�U�~���Qn���g�o��{�j��Q��r�01�{r�� $���M{P�k�!���wVLI��t�2W�)�k)�2G?wխ��"R�����|��� D�Kn��\'�M֐ad�q�V���ȃ�ˤ4�[��o��8�ڳm����E�Y�r�4~ϋ�8x�j��r|ĠN�:eVЩ>mY�~⃯�cW>o5v��j�����Q��;Z�b�B��-h��j�X�58�_�JYk�*s�J�ؒ���A��Yu c���sO���3��Z���9��yȀ�@87�W�Ii�_�m:1�2��ީ�#ٸ{؋�-sIM��>�<��zy��x�xfeUh�u�wLt1K��+WM��l*o�h�7�n����~�]�3(]K���>��5z�/0j�(�hG	E���,��#�)���U#Mbb�囡���4~��YK�w6����4j���Q����_���%�"m˘�}��m;���������+ʯ�(	'�e ѭ�PE�����V���Q�Jd����ź���C*�^O���>'��Kr��9��I���à!��V���3C��UH���fVr �;�x�|yI�����.:)�� �Ϧ+���Y��3�2������F�k�5�\έ��׵b
Θ�e}��Z�<�N�I����X�R��%q�=c�bu��[��Ew�a�8��~J?�Oj2	�D����htwĺ6Y&AY/���OFq*�z$UT�`��p�/y����]J_��xs(��B<5SB��I�:GDoH̒!A4�]�4h]Le8��Gz'K�h���8�`
��}����a��LV�yI��S+�O�_��L����CH&�9Vlg�R����׸�!��c��V�\b�轢��|��1oО�jvm���׌jQH��5�W���,ǩ�!��C
;� ��������+c��z&OD�-��%�бpS/�gpG�-� Z'�O��@M���u���b�pf���W�&l.7�"��F�{0��6v��f)_�����!��B�L��3��d�tab�S��B'��4����qn�r�x�(�ME��&@y�t�(�#\����O3���:���ۻ4��C)
yF��8�<?�m���ZJ�� g��jql s�u��u:P�V~+��C28��{l�#b��|V��K,є�b
�;��g�A�UW�<^_���dhk�����$��[��7�>�n�z,D{x�x��EL
�]�z]�<r��g�J�HX����]�ᩡ�o&khX��WHj���Ƚ�U�ޤ�����y[�KS��c���N��n���vm���g�ATe ջ;�h�����R�������"�H~�:������}��j����0���M��]���-N���XrM�7'�mjK.��<�%��[':���׬�]7G7�qےA2��u4/�mtnX[�C/��R�H5$I�N���&���<�:M��7�tm��h��(FBs|���Hєy۫s��ۼ�>��1:X���e�4W��)`��A�H���Z7#�S��۩���f7k�����k2}n�� �;���(��&������(te[59Y�J/TR��8��t߃1B�|T������V8e��E*G�i�tC�� �8\O�J�'�����E��셜	�'F�ˍ�]cr}�v�"t+| l8�H��!Wfp����_Z��.s�^X�	|U�;lWg��[�����t
�Σ0W�޴
��ӻ�J�����ZP�\�����ݼg\������i�>-������w�|AB%�?\\sY|i��c|���5Gnah7���ʌ�*l��-#4�H*gD�.�����BF�_�J�%��HW*7&�(�R�>2wG2��hN�i.+�$�T�:���^+L.X�U��z��80�_��~s.���m��\\�z5�e�^�Ԍ	?�p�U׽W �	�*VCz����÷�6jgi&ȯB�dW�9z&�M�v�6~��c=��9N������#��������S�>&D�<�=i�&&b�.V|�)��(�yK����[�zo��3d���''ӯ�K!���_�u���l?L�?!e��B;_��鳑]vr�W�xL��PV�����s<bA���aǏLH�qmqݔd�`�/����t=#���}�&�����L�+�?�65V��w3|�՟7�����01��N�Gm����	����&F6QLE|�ep��+�:!����`�"O�;��} e�dbG@d�r���lgZ���AW�
"�JBJu����dL���
z��p��12�g{mE��ޯ�){�:�ܘ㷬g�ŧy�."��:�T����޽8ۻ���LhZL�Z�
�Cu(|�� |w���*����8�B�|�� ���=��f�|���н��ki�/[�8Ļ"�X���>�Z��1و�7� 57fH�O&bE�'�_��#�"S,��2~@��[*b:�KA/8Is��_�ȞD��m;ѐ B[�9��NR�;ARm���w�A�{��%È�Iz�٣2�V���̒��b�:@��ޭAm�j��0���ʛ�U�/�B7��ց���)��3{B��i��'P�HY��KN�����D�ߕ$6�MU��X{���ۯ�,鲛
�����_>e>��R�.[��x��|ٸe"+�ccw��
/�M7�L1rmyd4��4�0�hi�IEŕ2I�`ˉD�|g�6L��]c�d�!ywp�[�$����F�b�����-���GG�Oᰫ[$Gj���
�q8V��G��zDZ�Ul ��`�㢔3����a9�?@�@���ͤ>�UݟB�G1���j�K�W�+�������w�k�ß����av�V<���'�t.D^(L���i
�b��V�b
��kfvM\9���x����?[,IG�7��V��A�=����H�L�|T���iw
¨)��&�eh�Y��;�� ����I`h�������A��$e3_�-Q����޴�i��+�2O�!���/�������C��ɂ]�砟5� �!��yZ6�2
q]�zK*鵇m��
�������2�L�Ł�`;Y��5�,a��ݻM�r1��D���=�HiN׫	�
�2�k.�{b�	�6h��>!��W<�̩�$��u0�'�\�]1�>��K,��ך
C�
M-P��������9��ǫQ���D���$� �Â��ÙA���:�]���̐�U�
����0z۩�n��%R�j��|ܘ����j-�Es#M��V~@�˻g�����\|R�b�xBţ�=T���a#� fehs��)���uBẛ��NS;��e��|�4}�*�w3kt�4`YB��a�s�X�24ཞ#Q��h�D�脒cB�g�<��Ùh�o�<1��'uC՞x�&��eF��ζN���'�*��wQtUh
s��D�]47D���J6,s�#t��lQ�q�lLI�%|8&Q�����X��N �!�s�	���+ib�^�O��s��X;7b��D��m�n.65��:�T�a��Ԯ_����a��Ī�BY�#���e���f�y��i�Q|���*� ����b�%���p�ؗ�����|�S���f�r�{�f2�
kb M܈l|�����u��e��S�i;�6�G�\_'Fn|3�?�|q��@�;W�V�9w:sX�����A�!�(���������eB>D�����vC�8ԏ���=�\ӫ���rB=�;���^�c��h\���}��V>�"3����h���&�i��n>����2������	���(,��i7"�Y��/Jd�ke�M��!t�3�T�Ϟ�M�K^�'G��o��>bL���FXw�W*���6�c�ܫ#U�Z�����M��g��7�Y�$;���Q�̓�N�Gw8Ntߨ9H�{a 򎰙t~=F�ԯ:w�G��LO�L�vRz-���d%��8H�Ӑl�ۚ� ����; 5P�/�LF�1u-� ��J@:=����M��a� PCoP�\9���{�X;�q,�ʅ��*�4�,��:B���;�.	��!�1���&�0?��� �M�T:b���K
�k&<�w�U���d����G����zS���n���Tb�%@��'��;W^_�����[Tx_�ڜ��}T�X����w1;���d�9}~�a��F݀��-��6%u5�ʍ6�pp��}5�|̈́J��'bj�h�t"U��k<��޺P����S1�V��xr
GxZpu�\4�vX�/�'���J44�;�J��!t���ba>X�{�޿'d�N(k^}�ר�H��w8����Z]�Sv��_���'��H���oμ ���]�lq�U97���9��E���~�Dԏ�@��{id?bx��P9 T��lƈ+��_�|����^�� '5�{)�$�3뷗S�w��=w^�;p9���D�,�H������8��_�uv�"���~���ЈI��yyȻJ��4�ښe0���-�:�i8P�U��	e�����%|ڙ�@;�<l0���r3�5S!<M���4�+.�&�4�.#x ��Ţ�X���pѵ���R�^���=��WRBM��ö�&J���
�FF��5?J��PU�*T`��� ��̵�1{�\��NJ�ܳ�<|�S�	��x�k�%�7@x��*>k7P�]3�?**��PDy2���S`��l����*xhl����ك!X��c��cE�t��+Y0�7�^��e�K�<�?��;m��!�����O�/�G�ě����K���W���(^]��m��ݮ.���C*�ym��)���$��!�i;�d:�4�1Z����W�W\g�P����N|U��+�+P����3�E��Ǎ!��ˀ�ʼ)q���$�3�!Q$v���A�x?�y%��?@�XòI��m�054[�	�-i)���$�E0W6e}��N�-�G�v֭�]Ax6j������ uꪫO�W����X�����C�C�!�y��O-���.f�i����*�˹,�=�Qsr�e���e��eG�}LN(�&�С���Fƅ% Ͷ�A��x�+r�W�0�`����p��d�/�>��1C�e��ܜ�#q�n_bH G5�!�'�"�9 R�,e��c7��	N��K�A�Zd{�FX�-�DtH'R�Fٙx�^����;���+�4belm86OU�[9]�м����S��W�e��l��~�B�)���l��,������ ���_�d��̱{w�W�*�ua�|�9�J��7 �?�ܶ������ȸ- ����"��r��D|z��5��³�u�����-�R/���FC4gsw�'��q���)v��'��b� �tn]I�囹��
�4k*"��>�hy9���5C��F�ARv@{�� �y�o�TR�0�&x"����?�"��63��O�T޶��i.����xM�F�8!��Z�D�	m٩Zud�itp��.O1�IC*�1j(�g�"�"�����8P�tИ���	)|.1K��;�_6.Μ@���_�XD"=~w����[(ۃ(��*��ь�CS8
�ο@����阤R�l;nDv���-�'1�	���0QE��H�߫��O�7�1E��$�s�ĎU�v�b�^֦X�}��w��*���]ͳZ�>U�ifƧ޿^�3O�0�O�c�60J�O�N������V���;�3k���$+�Zfx�1磸�_b,�9if��m_1.q�#���oz��W�6��7^� �V�tlg�N�N|�6 �qx}V�9�c�S�B�2w@�1�м*�M�����s���U�]o��9��� �����ܞR䗡(���_�篿��@'�/a��W�E[J�L�pA"�i�V6�Q�AJw�Oxi��@��M\��?���^�K.��g``��?):݂U�ط1Whꅵ�>j��8x���_��wAw$�9����s[!Lg>6zT��V���w��q
�N�	��(C%��ON�Y���"R�U_Ba�`�K��v�#���	�Ԑ�oq%�4x�b[�5}��D.���A�ɋ.+��շ�?��<�.��`��\�E\�v�ɭ��ޓ�}z"ܯ�ŭ">;u�ٴ���3gԔ&��c^�bSrz#�>���Ϙ����vl8��$���',�e͎$3V���
Zv����*�#P���3���ҧ���� �ycT�OOy�"L��cY�.W�>YxX=����)��A^R'M��:�Z��"���Dd�z�/��Q�s�?,��"�����{�\�=	Ѩ<�#ɰW�h6�N�t�3�H�6
� �G��/�%�yi�&b����L�����*�QۗɨW���S�nZ�����+c�&���C��;{�洄�z�6�\R����Z�C�OM^�l��T���>h]oꤟh�{%jh9%|r��)'�֡�hQZ���7�9aS��]�/���Ah~ �/:y��u9�h�<�Z�l�Ǽ��eP,����M���'�%�p����=ѧ�;>�;�P���{"��:�ԍ��$��^��YHjf
-���;�#Mz&�l�ǁy�Ȗ��G�|=Qۺ�Z=����+|?��Λ�h�����/%37��y�&����%���'此B6C�b����C��?`�o1B�����D�b�F�M�-�'=d��Du��P(mQ�x��P�?�qp8Qo.� ��PH�G�'��t�����v���}��̲�9��9�]U��րw��a�2/�	b�3R5��}Ќ��ן5��ؾ�T�Wb��#J㐩x�U%�J�IZ7o}�|�U|v}�'�2�a�����?C0%��w#�+�n�悲�i)�M�}�AXPc��r���`?;b�!D�V靇5�Mu���M���LwI�͎�2�Pn�6�X����MJw��V��p��Z�,�F'� a�{+_Y�[L��S��O�-�?��{)�Ꮛ�`�O��N�B���f�N���G�	0'>�'O���Hѹ��k�zR�Jc� Bd��pV�m��K�,5����d���b�ڹ9��d�Wg�O��R �
��<���r���\���i�����E��`Q(��<SN��Bh�	C䝷��N�R�_��@
S�f��1��ͮ�|p7�u92�����D{�g��6�'ٙM��iv#k�{{ڝ���%>�*��Q�����JTMƇ��� ��� �|U�U�d����+�A;�C��r��(H H�+\�{���/jYP�d��#��a���-�ޚ]�t<>r/C�⧹�C����uwO=XF�nP1�qb�UGU�iq4��֋(pM,����$;'],���K����nD\�!�h�+}`',%�G���8���ʛ5�$l��Сzʬ."�����9��Yqh_���p�iv"�x�ڽ�"�/Ƙ7�f�Ƶ�-�J������"����l1��%z�f
%m	ɺ�E�������tE8�	/3/$��Z5����tYԥ�_�-6�Pl1!����2�0�"_���MCJ�,�"� �5����V�a���y
���a]��Pj�{&�;���(�J�E^�
+�%-��0�JbLi���������~�8z2�|��6ʲ��f����nY��/}��O9�N�;7q7K� �f����� \�x�a���й����c3U�=�_J��=_>RoK.�K����3٦���4�(J���i�!�+y}t�PH�W��(�+n��X�#�ݶSj�"1�1h$g1R���bŧ�Ol���_<s-��N��`#�2���� �	g��`}>�5�l�W�޾�ANLsā9�8����C�|ɗc�	d�#�`T}����H�'�Ua<ɂ(N�m6�c���֘��|[P�&��������Z�ꏧw|p��@u�ʚ�i��P�u~���R�֣x�� nUn�Lu;�)U$�AG�����W��oia'����y�}�D��J���:ܛ�*��~lK����pO[�pj���v9wU�'Sq������l�6j���ZUqN0 S�4o^�M�ߘ����X��z�|�7&a�c�k�kku��h��ME�uK�������9�	�h�C��J~�~T�s�P�<P�h�7�	�5��5��Fk�1�bF�A�hV�7J��Iӂ6t�Q���Cg�~`_���_(
�x��Bi`�x����p��k;�_e��8��x���yE`s��(��xd�ڢA�L��

��p$���B&������Ϡ�0<#���$^gH��T`��y���Bޘwݺ��
M�<]{������Eh��;�\��Nћy�AD��,f9uhxD�
F��};����O�C%G�az�`�y+c`�h���=`��~�J�)�E�k �3�����_&��!le&#`�Ե7F�!P��%��?�\$a�Æ]���ͨ�
Yh�А.|oq�8P%,��"U�%��]!�S4�R��IqW�_��EV��Þ�;3l�S¤��Tty|�+��h��F��9��㑧�%��j
P j̐���Q/ƌa1'�4�T&6��4Q}�MB?�����ek��bG22w�)����1��
�	k��^?��~X�f�rA�&��{ӬO4�7-��.�)��IJ��b���� _�=4SŐ����L�תI���čgi�L��G9W�ϗ��6�Q"L!b����F��Q4�\���+��сmB}��0�Ez��I��I�@�w�(/��cڏ&�j��G�Ӝ��J������o����kksZ����厲�{�4x�=[u��8�pW��m<�� ��B ;Nw�+��)9B/b0b��)N���Zy�m{�k>E�����	ٶ��RN�Q0�P��0j~�O�����)Ι塝C�ϫ%����t0(Cfڡu�*��}K#�p�/�w�W�m�t��;)e3�VSs��_������ڼ�k=Uή�����$�E�Q�Jҡ
$�V��E�0����f���V=�1q���b-�~�[������j�8b(�֍��@+����I%�]t3��g�����z�Nr��ZR��N�it�.����qo���P�)�=�A�����/s�8�"k
S�!�cAYx�1͈1�l+�l=л��s�O��)��S���$?��K�-[F�!��76��$9R�o�sRk=�RA��iڽ��4w�%Q	�Lo���kq�a�h����J�gvĠ��8T�ǃ9_��9�����d:���0�����O��|.8�k>�$�Ye��(v`�
!�Q�Q���v�S��q�7n}f��� ���c��z�]Bݹ�+5��b%���z�y-�T��q�B���Ç�(�ɕ�ٶ�k�0B��mO�P�F��y*��^)1�G1���6��V� y]��u�B���)%��	x��IhrY����E-�~�z��id|�yqd���v�kl?����8Ĳ׼�l������B	��x�'�m���2�^pU꩚��h�T��>e�����j��i�7\?��K��/[_�����GZ��SwZ����|^��`�>,\6�ָ�M:����e6.QРƮd��.2��3���cޞ����	ȃ���P0@p�ʋQ`�Z@)-����*H��R<�x�e�HS�w����%�ŉ�M1��0<q<g�K�Ag<7���r]� N��O6�(�1������/�f��1��u�{8=j~K��X�����D�����/4r �_W"7�ا��-?,�T׍ъ��>�/��3�B1h����pYhh@����Z�C�1u,;���@����N4�1v��*���?�Y��X��`�}����D;�[��iWI�٭j'��JF�4R�������(�����:�6b�>��C���v^����>P=�cЇVe2�~S�(s�$pe�q�4>K�hq4y����uа�n��^��,���oӉ�r���/)M����b��α���X%�2�K��\�3�?��=��_��Tp��d�\J��/�罆��$��V�L&(lJ�m�i�;hO�{`�>T�Fx޺_�2��~^93�;�uo���m�.��I��P�%��0q��a�L����雒���mte�T�e1�Y�} d����G.b+��,��e��vYTP���m]~|(iQ�$XTWbB2[��m��E��� ��~%u؎���4K�g�İ�Ƃ��S�F��I��A�D�/�݉(�| ~[ϊ���R�ȗ�����v��H�.c��OU�D��[��4
Us�F��Lw��|uj!��%j܌Ʌ�9��n�a�K���ȇ���y��ӭ/3�E�k�s�mVq���E�ڂ���	J���IBrF�--k�'�����J��1�����tw{j�~K���o�Y�wy3��܀$+���8K�:_����	-uL��}�{���$��TE�n��}r�V7�� )��wV�\Xv�>;�j���S��IR��n�������wR�0�S�)ʒ��>`>zo�����v"�W��f�|������T�e|��u���|���YP�gņ��[l,���F��jM�Fy9v�Yx�gb��U�w�f`��؍�2���v촂������>jѪ�6�՟��,�&yB3��d��y�y�/`�Q_��!
�}�5f�9��7�{�;V�����eR�g������d���.@�GCÎyjx�)H)0��d��'��h��ܡzrx�2�����vTT�!D��R��Jp�eP�Z����;��0ߘ��b<`�k���$��Ǚ�e�5�^�f�Pų���u��m����r�- |����?y���mgF�`"�\�3(Ȫ+�Z.O��V��*�3W�o�����Wnr��]CO��$�m�����j��P����|`�kC���	�Q�]�I��k���I�wJ�x��t��_�]C��&BJ4�w�}����a�bٟ^vOX�g����o��Ǩ:J�Zd[#�䙄ߘ�U
�~���	�U����>��Z��.�}���.MM����8�8�D>>��,o7��`�;0ً?|��~��&�C)�⯜�������䖕�B��-z�!�r��Ʌ �����4Л??'U�����'��y����ci�C6�S�C>�k�ʛ�bdb��C.,�E�6M�L���K?_q�^;9ǂz=/�E���od��z "s��q���ܫ���$�� ��#��L'��'6S�i�̇K�V���)��1��6�j���a|���z�����7>(:�&`o�z�g$2�HϹy��82/�{/E1f]C���8�9�9���+A.�V�M�*��Q{'c�,����\���w�7���s������U�J�\E����؋=uq+՟��h/c��mX�.��QBM����?z��q�C�"ݦ&h�,#X�j�:�Rw�Q��L7e�/���Bs�������L����J��$VN���
Tw㷆l�xg���j�6 ���~ ���]� ��9�V�.}6r��0�R��N����㱫�9��-&������
bG�A�c,�
���>*��%� �f.�?���8���aj79�r�����d7Ȁ�t
c��D�A������aJ�̄��6��&V&V?7�����nw�eL�k�r��B�NrC,\��ؕ���[�&�J9���ƿ�^'�7*�ʝeg�@8:�%�H}̊�^�CJ�gG�A�0y�S��xn*���'5�.�Ҟ �(�3���X��R�0y��(��6�BR������ġ��t�֚��u�IT�%9�N�i"�<9#��G�u�-���d��oI$�HW�Ш�r���i����4�6n���~�]6���{�n'��u�t2�.5(W�{lܑw桫���b���WP:�,h��:��R��S�F�xZ_����#.Z�:ә��$��@�6�F��t�X=q�7d�9�יz��
Oq!)S�.������EΘ{�x�9����^�ͅ�JN#��"���>,�>�T�}g¨w�������ml	���g��^� �S��N,*y����P���� ��a�#�8Ek��j�a�'?刃�Ԙµ]����L+��n厏 �����S�c�:%�DQ����(�>,����C����ĉ#"3`�Y�y�ɲE�Z؀|z1I-+�6�h�5/�A\t�@ �t~�7�x�z"��%�m$!<R��A�Ƹ�Q2\�HS�@]��(z��=�=����>|�˔��h�j;�I��sk�1��nk�6����p*�F��,����HV�S��d����s��*�D@C	�7*����Vy)�,8lW��J�ϠGLv����e<�X^�*�#1�ջ��y��r��]��ɍ1>l1d�:;[�����,�B�7�7'k�/+aL���ƨ����
�����;����w��4pw�AĆI�q����۫��!��b1%~����wX�P*,H-s�Y�LH�/��E���P�CD��~�/"<
s���5�vRD>�����h�ê�1u,ҧ� �Zˎ�I��"42���,9Pr@�P�֓Rw`�&�',Q�+�um��0�z�Z�F��&��4�FDc��`X��<.���y �Y���|C�
�$�z�s����
�}<h�B�H�B3�IA��bd=���μ7�U�e2������f��2��6���wgV=�*)ݛ N���0�W�9'�iߋ|4���Tr1�8�	@��, �R�qE�=�eYøn`Vj���� ��9�=ٛ�a�w�\�D|rYx�~^��.�:�-�_�O�Mp7�K?N|}���6�2[{�nP�h �%(;h�Z��uy����R�)���d�|���2R�A�{����)�^���-�a�)h�oh��/��]���d+40�|{W�Ң(cE��Kj[ F��j�~�q�B�����s���'}�V��md'��D�vQ�b"��V�h�����~U���p�����6.�ʝ*�~�����8c0���D$�0��f����i[C/����ZYm��jڂ�ik<H�~h�t���#&�},v��SѲn	�s�}��D��X����,�[�߷����'��T����)9."�|AҎws:^�F����D�םԬ,~��'@��=��#��h�A͒2舐��-��P�~ĕk�5���)����c{w���~ڬ:�jp���Z̡�Ÿ��t�|A�%ӧ*�u�S��|�?�19�V���G0������_L����O�pC_�*��M"� ��35h��׻z�R7jϓτ�Y�!�އe߬��p3�6[�Ei����D(þ^(�S����x���-�&ʹ�M�#u�}��g`P�|�ʦ:�%  eҝ�T���c.�D���N8|��0{�;�"�v|X19!!o�D:(~:XH�ǧ�%lB|��k�Iq�BN��a��L� =8�}+�H����i��s�@a�5�	RΩv���u�4�����|���,$F���~�!bWB����d�����������C�[NЮ��pߪX,s���lA�x��ޕ>z���Y.OV���Y@2�����wv�`B,s�U�aG�%��TMߠ��ք����=�GU�y2���%߹_�|�����q�͎���`o*�����t:vD\���T
��yp0vE�AP���3��ƒ�g*�� '�9_����~�Ɏ͞V�c}*Ť�W83@(m#��&���NWŗ٨s!m�Ǭ���i��v1�T`���q�m��9��WᷗL��՘܅GB�-y�����I3�g���\��G5�V��YY �
+�SȂ�}y�޹�(�I�c�V:f,�VU/�������`�� t����#c��r2�5I��8���+��=�,��6u�!J�A�ޒ��J�;��/:u��겴,���1�Hr^��^��W�/ j��_|$��xsT�J�_ٻM�@i��Ia�0uw��"�}"���!�k5���z�Č*ƒ_�ipD���垌�f��.��P�y/��Z�Bǡ��UI� B�v�\Ze�i5b:P�E��
(��Aդ�����{C��X�����w�j�W����T�u�]�@+�a`�͖�����&#4�)��3�Bf��ԯ�Yb�~e�����Җ�c`��AЄ2$�=��x�DrJm'�|$�n�����ī��'ˁ�]OE+�o����X���*�C���&���Q������6M�}K�<;���`BS2�+��7@����+!�Vy��'���,F
ہY�޵�sR��
i���e���z�����g�`��x% +���:��v�q�N	Y���P������f+�S~����J���#�0��;;����$��)id�6��R��%Q��$�U�8��$�&���"o�;���`�B\v;OƐ$���eR����$Sԝw�X�}țBZ{��� ���`U�b�D>[�����T���	/h�%]�pVH??7pݨ��R�|�yp!U�s���s���Î~�q��Xh2b"�]��T��&�76T$M�8�h�Ǆ���|���(���|�u�P��|Y�j�u��f��"��ܕ�����2|G�W7�3��u�?��k$N�F���N-*���V����fm�w��)�����+�й�*H.�{�Ӝ��:�_��K\~����*t�Ӛ<S8㏸^S�:'��9�/ B��sёU�,`�"�N�I�B�|N�L2广�ڈ:���.&Nq�i�@wk�8��p��x���(_'�/+Ǜ7j%�D��`<}m��V�,:����~PE�u�ݾ�Yb[-ޑ-��/w2b57c3Mx�wY�(�&R�|&��m4�R��!��&�^�ϩ��9}�*����ȧ�;�I�Y	 ��_T���6o����OƝ)��sO�F�q��ŷM�a�b��<L��L�q�8Z�B����x��8�@=����+��l46lڨ��G�g�����:���>�z�4at�j�p
�����_s��[���̏��	�{�ܠF�X6�1��:�_I���G�U �ʐ�$�f��4+�P[r�V�v0�) ���S��~T�����_��H�iRj�Zڜ���X�\4��������u?���wRHKg�Gc�@���'���yR�(�P���&ą�3�[l�>�����ߐĪ����B	���bx{��Ь��,���Ok����Ҹ$1�#�OG[X����9�P#n�Eg/ Ë)D�����N�~�I-1yZ>��Jbd-�x
^�)Y�AX��W��!�� Ÿ��vE�E����7X���V>�e ���2]�x�0�ס'¡�yH.�}���$�� k�-�*�����>���S�6)c,Uܒ0�7����B0i�J���	ŽV}�mp@:�ƭ�F�s��1����^��0�����gC�!��x�p�]T��&5O�^��AxE��* ��������3Hk}���܈�)=47�~�_#>�u�*=N�;���8���� #���/bv�7A����0$$���k���[��������Z!U��G�O༁�2P���Z��W<�h�)�q_V6bR�� ��Hå���)�BM ��������u��e�C:��[����V��J�ٮ��W���Tط�
� �',npO+�hC�Tƚ�;B�
ى7�nD43�'i�a����9�i�e#�nNu�^��Ro�0~���|�����,�T{v$� b/���^o�_�p��ÛG�Z�̌�Dۙ(���P�1Ib^����=����c���'���I��EE��e��pq��;�2�=|�ē���!���j�w��,��BG|K������ Xz-��Phnxi��_-�]I�� j4�[�ຝ��v��������j��0�=_��Ւ����˽�!d���N��T�+���C�k�����H��G5!�o� ��@�J�4�N��~���d��*Y�qF,��M�y��g6��'�lS%c$k\p��P)�:m�(Te%�K���&\��um�}��l��[1��
I�9rKe��a|�O���wV1ݯa�7+�q�݈�C!��^�M?��<�
o��U�ު��+���[�+��"�O1�� HL�Ӎ�t]�Ե��X9K}�'�t��Y;�~O6���T�Q��]�p�9�<.��ѷHx�{q���vx�q�?��Ⱦ�4ga�`��L��؏��i�!�6|����y�g(�_1f�gAx��H��I[�Cn^ݝ'���r��H�FA�f��ijl��&U^Cѭ�h9�.�Bzk)��/n�E�z���ʸV@{��������g�(ZA8�?i�y�n3j�6I˘c�6π��=a�;f��=
�ʾ6�=T?K �����k�=B};��?"3��gL�S�s�U�-|�6�jy��u�7���p<_�������r,��]�ty��}z���浊�jJi���시hî��K�0��
K�.%a>E�,��K	�aAD������<['�Xj��`}6>2�*�d���l����!��ĝ�����;x�Ĕ<�i/�q ͒��AK*y����΀��|'�[I`��������"�CGjA��o��`C�łש��iS�\�՟���S}O6�5���*���d����/�������Ն�{�F/�M
^�����Qd�n$;P�2=�C@�U\q-O�=��2Hj�+�K�6�걭&	���ӈ&��<�~�yy��7�#��G.,b���F�!>s���8:m��ծ��+�>*�����Ʒ�Jj\^��E���C�Z]���uZj�m*�i� (��͙�(9���/p���%
r�F]�M|�]1enJ���;c<!ەˤ���D'T�7kkH��l3�}sO�ɤ`Ђ��bg��/[]r 2���\L��;Md�#����g�x�.��[!cT�#ܑ��.8�SA��d(�j�����x�����)5�3����4�9�k-壱)����h	���b�Vb�"'&!��C�N[F��:��Z:�x@�j�U�#�4�p!UP_�L�Q�� ���./b�,����NM�H(?����SP�>��+��,��q�;���s����U�[ϲ�'�Jq��ӵ"�r���¢�a����P�Dy���,z6�b�����kK��l7�R�S3�S��趆Aږ_4YV�)ժ���h���V��T
l��/�Lfט�*�I0<2�S�Ԭ��"7��2�u�:v%��%r#:�R�$�0���[����"��+���P�X��dq�1Y��@h2��O�#À����ӋDj�����w�
r�r�A���ؼ3]a�Lj��� ۍ�D���Oy7>�$��J\2���8��u��<2���n�5"��L,��$��� �ڒ{6ˠ��;7sI�|f��#>���y��a���f��i�;D���'ܺ�b��ЀVN�2I0J�����'��6����}�-Jh�ĸ�3(�׳��rZ����f�ń�Q٫,��a�ibЅg���������z��5(�?��!+à0�n��Cma5��ǋB���������z|8uF�����z7?s>)�Zfg@� ���Yr�X�籈*-���'���0�������*��ܷ��lP�o��a�$�u�PH;��0�@�+��[yWey�^ĒM�nU݌o��m�?sA{���Ak����/3dس5*Wq�k�S"~&c�,]`L�꾘�z�T�rK�lG�o'�e�p�#�	Q��~�=\��f{tj��-be<��2Z�7�vܙ�~"��o#�a�h��XN�>�n~IY���e��Y�U^X�0��k���:�~��-Q
G�TG�+կ�J�l�V�����|a��Y\[e�9:V<Y��եJuc����0����}��Ӈ�-���w��ʪ(=mM�X�����E�!��΍���S��4�HWgr<R`�.z��.���<�(����	j��I��0�W��u	�>�����2C�4%-sq<�:��4F��K���&3<�>��A��;B�6�mOq]0Ċ����;�0̈́L� �3�o�����6�'��j�v��J�eܛE�<zԬtQIN8i�3�c�Wҏ����`/Ҷw��R��\��W���:��)~��2SR����V!zg���;���3�=F�e0.?UcB>E8��O$���V�/h����Y�\�jAs�^�j������ �`�%z�D���MpK{�v�1u�9ɱ�.�.u���Y��� �|�����OPo�o�X���<!�Q���)..�z�}�e���P�����Nb�i��Gh5�('>�}Qb��//|�x�R1Ecl��!��~P*g�caKf��}.��Bh-�D�eehp�YY���ø��:Κ1�_(��v3����˱��q��:�-�4�#��ᘴLi���Om��w���v��ք��(,-9�t�I�R�l9���r4|�-�60��As\��p.�ɘxfc2����!X*I(e6��2+����G?�+`�KE�p! �-'9$�BnD��x�����ݸfW��w9�*<U��铖(�[���IAݼ'��mL%Mb����X�ׂ�	�c���nԔw��$�k��2��)�����|C`}�Ym�inЌ�J'�RG�S��i�����HRg�\�d����Y����Ǟ��]���\��������m8�ç�.4s�A[�3�T�dI낻-�/Â:���e�zj�[�^w�X31�g��pg�|�Q =R�u����
D�V�Hju����b����Y��f���IB��k�R����w�S&\�Y���;i�q�bAi�"�����y�%��G���"����9�����Y�5j�O���v�\�Ca�8ψ�&I�o �z���V�^���Mo���m���eIb����a�_E���=b%�Ɣ��+�^X��oL;�m�{&Ni;پ:}c�0�,_!�)#���_�I�q��_�SLg��lo ۑ�=�3u��w��i���3ԧ��6s�D����X���7��"n_�K;�!DXUH�^��8D�4;c,!��f"�]|i�/z��~i�~`�1�:y� �h���0�.��ٲ��h�~�M�����
*[p���;���O����崂1�=�5͛-�Z߻�����]�n�@@",4I�o|!L�9��q��?<[`b����m^U��E�Ko���� ڂ�U"�̙�c�����T�C���R5A[���@3S#�@R��V�t�����ods!��)e��wͥ)X.�Of���EB �㤉nɦ�[�̾�=9�+����t�Ѻ1�2�dr�<IE04��S&�ߛ�ĉ�_�S������)����$F�5�C5���:[����#b ��	؞J�F�r���0e�P2�?ON�v��t�����8�������_���
ЈMw��4�GBN�t0�25��Q##!+�˽ES�������k5�&E��z�HGR�Wǽ�ϣw�r��е��)Xn���ԛI�6��yp9a�U����[�U����t�x�`-m��j5ڌ�c�AVPo����Nm��t}ڧ���v�H�?GVֻ7�a����I�x��}��	?+h�i�HX��PE�Hg�#��~�l�xmɇ�e�v���D����))<�1V)��~�����a�Q�,�@�H���&u���j[NeH����/HsF|L9?g0�:v�Z��!,!�ڡ;��o\z[}���XOe�|���$&��X�QH0r�!_n
z��7�&vE�+��d�,��Ń��%ߝ9��gt�m������F���gG����ks��2�\�y�3|�b|�c�Z���3�� �M��q?X��9���/80�B��ȕ�{���mW[�}�Z@�H�ֵ��ň���$�Ȑ
�Ƣ������Wt�������s���6%�BP�^�qWwb���Bϭ7R�b��L$� 9RB:�9���N�*Y��Dߊ� `�U�ы8�!�#Gw��|D%)�_�0ݰ>��>�
�j�]R/����X3"�F�pe}�d����;��	�2`M��7���v���gs%K�A=צ
b�*z�ǎ�V�A�د�.r�;�E�J���%n��S�Q|/Ծ҇@6L~���3�<̑�;�ue'�s%g�F>N������r>
^?䢟���=��� �����k`�8���[�Bwµ�������j��ny\+\՚y�W����������,����X ��H�T�21���xQ0cj�;�{-���nmƗ۔VĩcN}zմ���|�M�/�yV�q��J	�BSX�5��ѷ�n�B���^�=YgS"�n�$��y����=��BT�`�ʀ ţo��]��M���R�+�.L=�6��!����R��Z��J	]ٱC�q�<�'���]��q��T�D����g^�:�ӊ��f2���/A6���f�>��9�׻�[�� H�����6�[�e"5=w�e���3rT�u)��n����R�t��A͓�
D	�������3GB�e@�K"�M�)���4�O�-ԠH�Q����VJC���"A뺬*#��fk�Ѧ���$�Rd���O(k1�4�߯�U��3��qu��MfLv��˧��'�2U�A�]H����{�	x��5�*@6y�g�
6
�H�4�����������T���Ud����y�A�w"U@ZѸ��0�H�i��f8G�m����f~��~PD��B��S�v��uR"%�4�%ug9޾6�$��y�p!���־�C5(��}��\��׮/�+�<G�[�lq��3&�Xhv����_�"���%�2�|1�K@�Dj�&�;#�j,$�HV��8��Y��-���q��3)ϤZ�I�����}G����-��'��;𠒰�UR�?��a�e6*�a���#1���d��u�����~�ס̅Pq>>�lx���w ���b���O��e-|؂;wGX��H��l�;ʮ��F(���Ь����z�:񹪪/a�1��ڗ��ƽēA��d��2}�7��VO3�mn���^}����b²���P�e�싞�ܟ_�n���+ ���>��m����V~(@����:� �?�/�+�FS���&��h,!��tg�%�A�]���.�*���ؿ	;�R7g˸ �OW.
m圅��ԉ�sf�,`m�Y�y�'�}p�����I��#Y���ƶA�x���#ƃt�Z��M���ne�E�$�j�8�*����X�V�wh��H��Uhkn�V���#���Ϟ�N""���=����o����]lRst��%�+�f=�� �QS.�w�~�Th�$�����Q���R�9�3����)��B+0E�m�ى��iC��l64�MgH7�Ǐ��\�m��r&wi7ɮ���.�m��A=x�O�VN?6�T<��W%Ŗ�~k��2�>��vH�u�Sã�J�&n�, &�Y1^զ�*����H�v'[!J���|�A���fω0����Kd�S�Zr+�����U�ft��'�V��U��jM�Z�K���FZ�~�E1�1����{�j�}�*A�J1J�ҹw.R� 5��wV�ơ�N���*_N���^�H@��ժ�)�����[�Ý����nj�0��m��d��2��s5C��w����iaHQ�V:h�\y�͍y��[ �&�������eT��E̷�0�(]O�W�������L���EFg#$B�D7���pKc���{����Q�����4�j�i�y=�@=Nj ��T8�Y�o\*�doy��{E���gf��߫h&�6]��'&�[��T����L�H[��*��~Щ� �>`�d_�y ���	
1#��
��qZl�'�_��s�Z��ݹ�E�UEgw�+��_�试$,W����b�F^.t@WU������6	x��l��?m�V��n�Bw�.���c��Q�*�y�d�.--��$n����Z����k#e}��Y������P{䒘��#���<�=e������?481u��^R�bM��l��5�k���fu�����o�ӌfj�I�,�]���~�0����J酛-�n!�v��pп��.$��A��ÙHM���801�TM'X��ze�.b&޸�_o�-�c���D�w�z�<t�����x���A]�ƙBj�9�a�˻�M���K�3I�����Q}���#������$��焄*v�P�4���(�q��ST�6p�{Zk�	��Q,m%�Y�= K���]�
,��qլO����P*�8��fՕ��o"!�D��F`C�2��a�����B�c~�E4Ŋ����8�e��D�<1��uDYhn�^[�Z�ǃi:z���K��}楽��� cA���+G���@��������/`�<lY�@�������qriIy���P�숖�Ex��y��$>hKpɴ����$]�<�֛�h��h%��`��L`x� �E]M��_�%��e��!��������*���ͤ�,�u���xw�zTq���@��S�mN�[Ʊ�̆�x�Pd��p[�
Ѝ�sP������Ѹ�KGLB����!�ז*�D�M��r��o��������4���e�W��X�=_/w&m�#g����0�ԃۦQ�,a�TM��j?�I5n����b}Kaɝ� 3�۷��aNx���vL�c�]P��?������W�T�H�b������w�k�����b���N����ev����whRU�ʝ����"i�_��{��sE�sB�'�RZ�Z9l	Y;e��q�BT��~�[����)���D�0yخ�B��Z����g�>e%��*���:v�&D����<3TCR��Z��]�ͬ)4`��]d��y���\���E��_��E�)i��̍�%�rC)k�@�t�S؀x}7��^��p�f,)F�yK�@��+�o��Uա���\�I8�`8�x8Q`07��8�_έA��J��+?r��(�4����Y�Ts[�OT�QO���,�w�����$,�4�>+��@���5�5�Y;8�,HӡtUW�����r���=�Eϭ���g�IbN
l�貑�{���$�t6P�:b3#�����ʊ�!��Ȃ.�:�?V2�m)!+�@r�����J� �⒠��Ց�B�g��!��>i��̹b�T���j"�%H�+ʚQl��[=/�.�c��7Z_���8܍��@��c����dɰ
1��~���3��ވ<\N�kb�[ӄH��o���dQ�
��y�?4ms�C�_׵0�)�3��{��A�(�2
R�X���n�f���謫Z�M�\�.u|Ƀ������V�Z�` H(IFq���Ax3��!Y�=O��D ��P�8��c���)#����dJ pR��\Ź2o�����cO�ޠ�81I�!ұb4�JH�M��$c/X-�i�f���¶o�`���9�%x�m�/⃄��x'��`R��F�q��n73��Gt��%����OY~u82�0�4���T1�5zz�6/�AƏ*����DQ�Nyk�1C�pgBf/8 ` ����I�Z@��=���V���%v�{����+�ЊFp���m4�i��������m�j̦A�����>����V컀(� '�v�UH�b�n�[���������z���z��e����?K���Ճgt�z%[�:ٚ�'DSt�پ*Q��=�],���8X�x����"r�
�6�H��U>n�"ڤ��,KY59W��;�=eA��/�0p	�ˑ����q� ���v5��}]_�N�:�	��"��&I�>��:I^�Q� �%���i�>� �1����wӼ�xH6�ߺ�	���j/��W1���-�b?��\����u/�9ER���K�i᝜��J��l�sv�\�=L]iD�/{���<��1ļk��<�8J>r�\Q�\�UUM0�@E����(�:4\��1���fV�d5K˛Ҋ�O�ՏsC�QLj�7HB=L!L��B��`��y�^��w'�Q�Ժb���8/��9�:c���Q�7�X�sT!�%6�c�.�]�4��M๲R�8:���ڐ|��V��bܵ�˵{��l���M:DP�G_��V�(�ط�s/������镖�^	y��(�^�+sh��_���\�yd\N�1?'�T)*%�Y�P �0R�$ U�ӭR+z����k�F�m�4UTE�B�UL`w�68ʏ�7���f�I�s��q���3�`�h�cb��ہSn�O$�X���*�����Φ�Ξ�=\�lwp����z���15�a��M���(�y�>�l�Ti#��$@�k=&6� {����=�L(d?H��	�����w<�V�͏ ��M>\�u�1o���d 'J!5(�9X	��u����,1{��n��c	i̙�+;�C�J(��5p��Z��J�滊~5�G�f���Ѹmn�<��c� �f���FA�a�o�K��uX�JMʊ�����}P-��?W`�k�aT�k,�iD �%=s���f�Tk1_)������8YI�'�Pi>�i��O��L��UZ�
���(��u�8�''=�
\�8�/C�����~7b���>�B����"��\q:B,@f�Vf�(�[Ǌ�D1�a�n_��3s`�7����ya�~Jjb���r{��s�)�D���%�.Μ%��y���*3f�h�Z�ݑZ�L�k�(��rj�hk�I6y��'���-��W���� �e�f���\�8V�?w%Z1lt�pXRr�i��{ÿ+x1A�TP�	��897=z������A��K�t�H��?m.�����5{��a"Lƣ����Cv�@5?����$`��y@�3s#�'JUc6�>�������߼�5��(x�Y�n$�:���s�BV@� ��u%��i���!�l4�1r�Y�f,��;�P<t~��ھ�����e4��O��]�gε�@Y4�[g�Y���@*=훻�*;&�Y������Kʕ�#&��h5 �=#�WfY}��V�� �/_!\E�7��~x1�(]���ފ���?i��'(��/� ׏|1� }�AY7�0>��ト��u��K���9T�r̩*��r���670s��s���L��A<|�25�=�����g��/������ا���Ӿ�!
tZզ�X��%́�X����[��F���s~���#���S�/f~��+�F���G29D���ߠ�X8��'I,{�wr�����k�N�Y/���^B��zh��y�C��qD\' ��J\�՜9��)�z�o�a�2K��a�~Ņ9�Uй�&O'�	5PjY���"lǓ��ր43�6Ttq�;uT7����i��ϊ�^H����4~�H;U"Yx��F�4�X� �)����5F���<j�ӻ��D��J�lT֖M����`l����sC�����$f:��<�;�J�	�{ˍ2%څb��=�{tG\j4�U���Þ��z��1�{�<�0�5�N�Wj �Ӆ��̨��T�t��|Fy���'S(�I�6�&s���l��C(��5����6Q�R
n�х\�iR��Y}��Reɏ�A�S|P�CHf#�wo�9wAJ����_.�/ml���0U�Z~&hY,N��ZJ@
:ݧe�H�7���`�La���i���'捶� RP�yd��V��N,�$(�n���6������t�X(s�o���J�A������rZ2��2��!̋r��D=6�*�{����aI2��&�g��ԛ t�9f���٠�4�w�8�ƾ�����"�$�9��y���+3���s��ͯ�\kY�%�Ԋ�1�SI!�S�Fr��::�Ł���@�.��ro1�5�'�S{�Х��"�	�8I���<mGȤ�,��g*^�=yWI��\�^?��V��5���&���Q��(n�e�H�k c�=��_�]����X��0��{��R:��TQ�_}����]��;C�c+�n���`m�i�û���085紱>1ĉT`�/��w��rJn*s���Zn�R)���ɹwN$�u�\kJt�!.&�����q���e*�����+�`7�6/�p������g2�
	(���T�	Nw���hԆ-�7(��x��L���}��Tφ�t��������i��#d�M&�O̐� ��fƴ��
e�-k��茿�źK��Ig��e�²�� F�w`A��
��n��!ݯ��<�d�{�!^z���%_:-�r�ɞ��̗*w�/Fp�%�v�q�Xi�/O��Zy�'�l�ҵN^D����3�S����>?���������t�Cv�������E�-��Ww��G�,Q&�j]:P� ��btr)��	ua/���A��K�'����x���c7%��`|]�ɶ�yrPP�/9��(���EnG�>[��
|��UT}:�X�f9Y���r���a}���ܝ2	?\/9�'���-O��@Pp��B�������$��x�I��So3�䶝3���V~.��)U:���6�����hKmB�ӆ������b{f�'`#H���{��M3���"QY�!eL	Ӛ�h~0�w��{��9D�ݠ���d�&�	�C��W�TTE�	�t�=
@�]t*q�B�X�%- h\-%
S�g�t�#�w�	�Qk2���.(O���ыejG��kK��p!o�Zc:Y�iP�d���H�?���r�[D 1(��ޣ�����M�(���*o	Iep6H-B8��獋L���<�Ry�57O�۶� 9�����wH%"-� tߊE��nIQ��-W�ou�).�Ph4���*��&$=��gtb1�.�l��Ya���҅�kQHOg'�'-H�����eڄz�n���f�y�9`�Ww�������M�%��4��H�Hh"��t��!�F�����5^�H�6�=�%9#Ŀ4���h���u�aT3��yS�֓.��w9u槊�)-�R��`����(k3�Sw8�͠�P]�'ɂCgc���)��f����:�D�B_��A9EQ'�W��%s:��}�勀���Ѱ��R�O�5�?Mn.��{�Cs�S�J��J������8����|;Y�D(�j66C�Bҵ��4��q�)�2�[yvA4�vj�*jЂ�{oY�ݸ���Nh��~y���UDi�4\e�i�=�x:��4�z�A���o_dL�YMnvo�rq5fH����ܶ�h$-��R�5�չ�;�?���_���͒B0>s���p寈p:��в%�^.���m�6�#qNy�s汀��$�}��;����;P�^��_�RǓ��53�E��],$��b_�,�)����e_��Y*U���1x7lΰ�+�?�r6p�Ŋ�MJ�X��O������L�&l�n���8�]����@i]�%�z�|���|���MȮ��$x���ðM��(��Ba�zvLǖ�LUq���/�� x�Y��0�S��u-P�u�|��iaeku�3L�S�H���ق����`�������Y~�Hx��x�j���oٙw�C����9ց�N����O�0��B_�H�.�h��I=��n@������}��Ƴ�R��%�r�%Q}� [��*Nx�@�U�H^`6���R̩��f���}�7N�cj�b���.�ڬ��7�|�~4���2�D&.�ΰk���D�@e��V .�����{#K��wWq@D�����r�-w�M�G*ۤs��6�`f��KV������A�1Sb__]�]���-~X�U#��%9Z?p���D.�BS�]���g��1��+#f�~��N=�U5OE��vOt��R���+(�� %���RT0�0����B�^�J��XN��n���t_��%h&�0�nB�R��b� �?,"�rz��p� ��r+e���9V�\!�WN�cO�Q!>Q���^�hS��f6��Q�����2�B۵�6�]�"VqۑM,%j8�f>/%�:-��|B8��Y��G��TY0�J�P�>��a�d�� nNtJ%�B8Eh`q�g�c����Kc��l	�yYk��~�Ö��f��(����|��j����s��s���1f\1b���٪��CH ��zk�{Z��q�>���#�w���x������A�
�^�CLė���U��a�RX{��u�_�4t�d�PS3/UY��L~WO*䟯��٪�ª'���z�>��!V�F��q��J_�Q
�� ��ǀ�4�ߐ�^�!�L>3/)S�}K6�$Yq�^�����C����Ҝk �p��z�rۏ=f�.�O�ٽ��f�\OC�Y|���p9�J�t.u��7�q*�m{�����/����z�BW��`�RU#[�A{)�.�vãbdزX�1�1#���~n~�I�.�@�-~9c���Y�\��!B��Pk1Ic��9p�G>������<�[n#�ps�rKb�u�a��W�/!�@1c��wũ;��&7�ObZ���]e�~U{������,'�r7q9�<�vհE]�KD.�
�ha��"�.����(7LJ�C1����BW�3Φ���%���!���Ϧ�n��^bU�j@�K=1�5#Cއ ����&������}>���~,Z>,��С)ܩ�6���^��v�-�&**ҽ��7���N Sܞ��+��xjn6�W���+N{�=|I���ׇ��{w�tPhB`5虽s��n�p��BT��f��1dK�&-W��G��U:���_t\m��� �sh0��x�lj��)M��K�=\���Ρ�	e��o�fH!��{�ٛ�/_��'�	6X���+���iA8��#g�o㶄J�$�T����S�i�wdZ��O���[���Rl?��o�W��	-�i|4C%��6��{U�Ӭ��fQ��n����?�YO�A���>W��=�#h���5��P��k/�R�rV1�2�7tګ!�`�7�}����S��(v7;R̠L/���#��2���߾&��;�mɒo>w�+�|6�|Jt<�;��ĕ>�<ji����rwǯ�[g��kQ�/Neސ�u�VK'W����k�� �V�­����z�I�FΧ<G��zå�i�t�Q0���h�P�l&d�>��GFy��Jf����[�C�Z���f���)F�'�����K�m|��9��]P�&ud��D��N��!�=�A��w9.�����������p�����%��!��$4d���t�s{k�	xp�J2���͡ϻK��P��m�Qtx)������* �2�Q�����vz��S�I.�a��<��U~�]���L�,[APtn�υ|�Oc�g���G�G�L,&��`����O/Yah���@����ܽh�h���_0s]�(g�?!""$�6����qz(xǳ~�wf��IA��Ij�b��=���oNK�AH�uU(z��%]Q���i /-�[�E�t�3Bj���f�a�׺ͻ�D~n ��i-0I&|�A�!$���T�' ���O����v_hЀ(�%y}�ʈ%���x�4,U��_��l�$��� #�C��/�_�F27n{����A��N���];7�;�i5Ҏ�p�򆴳Y�W���P
�v��^V����\x�yM���6m�ʐ"W;~YP�_{��^sg;�qAu3F"G��^k�������N���|p�+����`� gh!6�XF��Da�$�~�fT���5�쁁�M�-k�[)��"%�Jj�&4��MISB�m7rO���r��w�t�	�=@e�����Y��
�JC:��P�7%P���z�/;�2�y��7�A�b�a�[�bT'��6O�ʥ�@��^�p��O����E5?�B�i�����lM �nHY�P��
�5�׈�Ā��UJ3��{������H��7�3�)��H��A�^���i��ZWA��ŕ��Ф��%���-K2��2�	������m!��ؤ�˃>h_.�8ߖ�5	V| ��ht�8�y�`x;��=����$>5�J�ob��k���dTP����t�_U���DV���>Ñ�3�o1�;�o��m(aK������ʐV]g� ���{m��=�yE�}m�N��_5�q�ђ/���g3���鮛�1�{!��kE���I-��=7��KPJ�.�SV���oS\"���3���̴��sf�z<�p�����-n��slg7��T�ʪk�/���RMz�}5@F���W���a1�gbT�j� I����s�R?��ŮIg[%kM���E6���n�.��-�f{���gUX���9��UN�`$lC
���3H}�ꃖH�<ݿ/Z��������
��gF2�6b���hF�P������M�R.O��/��<fmk5J���Nz�[4�с؏�`:	_}	���S�v����I)��#s/4� M<�/dn�1$��B'gƏ���_����߿�F��J��<>I%c��?����/U�,<B�Ӗ�_�\
����X�5F�^�7O%*xɡ{��-q<��M�2��[�ri�}ݞ%�Q�N�يv3�L>�?��Q�!fX
��)�:�g��K�r:p�@8���:[.�\�C�ה��� �ZG���d 	̭AB�U�������Ԋx�!���fX�҅��c���P]=�ԋ���݃��] n��Ik�K8��u0&��6A��Ե�pXT#_7��4RC�v�׭�(7�ҊR��6��en���ɁA�&��}F��en�+��ƍS>
/|���8�n-5�m*���m�H	P��$_?DT�լ�%���7���!�G�����J��܍a\�7<�k������m{�9�����=��a h�k�b(2�鹻�0�T�9~Qð͜+6V5������*��2Y��&{�y�<1;��hT�x�WėzV6�|`HC}~�v��	��C�M���#sz��]���g�ˁ��b醋�2��(JWj�1�#k�A���	h!�&���`:^��Q�����7�f�(9�EmW�ų���O�~�

y�B�����G�R+*[�P� �:��}��g��St(��,���p�'������U0��e	���rA�u6,��,��#�����F��8L7�ec��ߋ>]��2ٔ	��;�bO�����igшT S
�o;�{vv�>�26���J��,C�G=�.����Q�ֿ
L`��s��A9�DF�]����,�:\�y�����e���Y���}����E �9���o�g���CyP�!�<KĖBT?v�3^@ea'Yku��
��"C�f'�r��Wx�9�b5]\{�XS(E�f�z���w�2��o�;����}�h�Pp��� 7m
��{B�`�(�~�e?� �.W!?>E�X�J+âUX���,{0`_����h�����(�Q<T��
�8h	���Wu��9|��Co8!j S����} U�oZ�O��)��7ce8\�"�I���}���>�~��	�p�}R`W��<4�>A�`�_�E��z���[�V�N$4�sɛ�o)Thl����aD�ڼ�ue�9�	�+ר�QqO�5屚1��ȺH��X	o�n1L����E0��:tc�@$S�OR%mc��r+U�Y�FCY�D�ǤGħ���Q.n#pb]�b�ˌ�(,����sè�I�D�r9�x�F�`R~j|Ɲ~�k���R�QZ�eP�:9������*Z rƂI���M�;���Q���Wp_�q���%=4W���u�'8���)��3���b'mS;�9$�'3��qI�+�>��'���(;&$#"*����5'�ߔƗ���OũT!�bH���$��[�y�ge���FeL��R������Mz�{53��Y�(�(Nx"��zQ�����_0׾�C��\m�d~s�u�=��l,���X�����fhL�w��(8m�1?w����x�H�D$RɏC��x�C�>�L��C��I\�}��s{x��0���C��,U<�F�+~P��ړe	�0�W~�C���BJr�e��t%^��t6&�[���0N�ҕ�Q�����9-gh�2Y÷��-WW��2Ϸ(&c�|�ǒ�s �v�>֯�W1��&��ԩwm�8������N�|��aYLG��$�G�5di�G�$D�_���12PJKGL)�Q�Y��Fq�ǀ�t���z��F�)�82P@%�_�(޻���g5�|���v�ݤ���ڙ�r��&�ʋ�h�C��>�4H�?�!���h��)�V1��H�t%^8��H�,����VCi�`S�O���-�
�o�[����g"��Vq	�	�W0߈�Z��f�e�D��� C�zS��;�jaKgC��[Z]۱(w���B~۝GV{�y���U� �`���1��RA�E�ԩ�>0�2b��L||�5�"���ٷ�
J'4�,zJ��!����g�E|O���7jɊ7�e5s��N�{>�OӼ��d`M�TK�Ο.��@�{��F��'O�}�ک�2��\0����8|1��C9j�Ӄ�`}i}���EfQ�J��H��DV���x���<��d8��,S�h�1�#����Q�	�:[U����BQ�s,��B�����i��#����p6�n<Wcx���wqD�o�9���C�y����O>Vb�GT�dO�Î��5��H4��6>����sb<���	0(�n|�`�w�P�b�O�З�D<���|x�Ծzn��#��UM؝)z����!��n�D(�t�s�0�ãS�F�j��e&�^�p� ۱�v�q@UdBg��'t��u��<�ά�E~��N�w�$��.\����j��4V�J���7�./�RL�m|�ذ�L�}_�O��[�_L��7	�r(�DAX�lR��> "����f�'|�6>}ƽ���1p��` �V�ILT�)a�y2��F9�R!#
�CL�͎T�A�{꫽��*�p�U$��H��+���1_%Q�AU�F$hubu2�H?|�O�d9T�(�f�3F��}�>k��<4�8׿�A�j'������4��tEP���Z�%`�sb��/���d��4��H\�}J�K��S�����P(�|%���bo}���x�fn�>&,�Ș{-\i�@4kk�� sz�XO�)�����_�A)�ps�x�Z���wnB��$k@=�,�D�N�Sv��>��q���rT'*�	�ނ]6�#����V�.N�1U4%%��Ō�Dɖ�y���Q�����k���D	s*��=آ�?:3{`�вB�zeV�S��꼝֮^so��#ZӁ���9Ó����[�u>G�>�?�^����>ilm�Te7G�UW��b�)q &t�֫�#-��௛�'\%��uE���ϒ9�ࠡW�Kט���ı
̴-�o����P4幰p�8�L�u�0��˷gy%$+D=`��2Ω=�_j��Z9��
��%-�-L-�ֹo��/p�!e��y�'�}��/>Nj(g�Ӷ��*f�&�p�'�4���k�Liz[���N���&�>&`u�'�"���伸l��S/�@Xz���ՙ�4��bw���F�"7��G�+�B�FBxԕ�5�M�tc��go��{�'���7�+u;\�^=�`����v~FGP���\yؖ�'�%u���j�J�Q:g��i��x�Åyf�R�-�����ī����1V`B��j���Q�&��͌(�x_�%��)4Ӡ��Q�0�gyb��Y��&�j��w+p�� 0z-��8l$nu�TٲutΑ��!�@�����Җ�c�������T�2y��(����aKy
����`��P��p��Q���O���bQ�ْ�佷P��5�Q�#�/�����b7�@��*�l~��a@.W	�i�2�ό��_!,".-�f��p�J2Dl�0~�A��_��a<���nF�
ڝ�ިc��N^2jྕ�N�1�������c�s�^���LLݷ�_p|�F��m]�)*��|��y�rc�jvS�jy����_eRM��̎�L dwq���_��iA��}`���"��@�hۻ`ڗ�R1���̃��}2^�i�ųi7W�}T���<˚ҳ3����������4�!(�3ƨ8���&�EN��ӛ��yh-cF��w���������"E��s�1/-:a0�"���=e�:E�zc/@�&u�W�F�L���f��=�m�T��7�7���)�4\w/�����r�&s&�:�N��Kf����������ur�j��.���������_1ؿ�������"{SD:#���k�3J�5I�����M�${��m�p�Ly��b�i�:�G4�ف�6UP-�����Wk8��R�e$�Fbi
�y����� �ѓ�����W'ġ�e��g�apFIE�Y���G�|+�ɗr����Oq�Ƚ�8�폜�P���������3��Ù�W�r؍w2՞̘����Ne�h�I	h��R��2�%_�y���
vx�~�}A��d�v~�VYev��� �j_���*���В(�Xsf#������J} YRj�y�X�:l��`�0
:�y��>pl �u�nd �-�*�1)]��vZ0��&������n���1#kP�pO��F�f�"t�ݮ�������<�U�i�z�y�-�������qx��|X�A�+K/���}˳_7������&H�.�����:	�y��)D6���@Eo���M��q^�ֆ�À�,i=.��%��e1ʸݽQ	bp�O�q�S�^Oɼ�eŞ��b�8�nG?�lJM�>˺����
���������x8�.��8n���U���p{\�f�%�1<#u��$�Z$�Vj�B/lC���b��5uNw�){�D�H�<�R���"�`��ix�$��K4?-P6H^�/:`|�1n�
�
����bh�}�.j�����$F�i� GXr��~w�.�U3&'��(@ż��Y�=����d�g���d�*/��/R#O��ê��ف>�Ӟxh�U���^)�B�O0��`��|�P8~���ؽ�\F�+)%�d'	�I7��Yf�^}����P+W�ӏ�MՉ( j3����$�H�d�~�C��$䙶�׺nb�/�V�{Ȓ�0��z��C@����7�v����ɡ����4��2��䤦,�������p(8(�]�B�l�Pu��e6]��ҫ��)	I�G{���q!	��!L@y2'z�6 ��,���r���WN'��E�H{(�Z���d��i,h�нI�<�L��X\٬:�ySJп4��=/��Ɲ�8������D��<�E2��i����^�d3*�YWݰK����X�U+0> �u%�F��<�ɵ��d.�{G�a%�8:��(��]���F�13���G�wrĒ�(j>!p�
L�C��A��gr����� �h�is1vF��vX��.?G��&`K����;~H��~������/��_e�
dc3P�a�M���/{�D�lѷ���zʿтV�x�9�&yv�+<Y��ߟ�އy�RI���I���Q]�ZE�=q���O@��^'Ɲ��ZEdV�X)��,}`�͠�9��(�!B���M�9�%'�<���;�Q��=r���V�^�(h���g��[���&�^��������G���kwz_�mw�++g`�w���D�n�]@�Q�N)��������~;�:���܁-X�u_������������&/BI*����<Gӎ4���[��Y�L$tc � ���
�Y\��$ˎ��&�TrZ�|�G��$��� b��J�0ذ�*3"Zk�����K#n�X�F�������
��v��#�S���rS*�=[�@p 	+��։��Ӆ�1! g�n���t�e�x ��}�{(��b2rhW���&���^ӛ�aL�Q�^����8bn�T����!�{a�?TW�L`!2�e�t�8�eZ�M����?��~ZTp�]4�\%���s+��Ddl;9�&͘Y�P��������Q����V���������A������Tu�v�U�4a�V�����W��O�A�ŎC�^��(���⥸�.X�
�u�zl)�JA�
��%�sZ�~nD�~�Ka�>]u��xp�Y�u�c��h������q�j�}2?�ta�<�vp�����T�kAۇ^���@s�h�>��(@�S1�m��/��
�e�\�0G.K�<"
nj�q"I(�G5M�̙��W"�Ocz�dM*�^��;:^;W��&/�H)��̖�RNNS�CL]PPO�r^�T}��0'4W�������'�����D�Os�X�KYV���Bg �Zqé83A�I̯-��	�w��E=}��8LP�*�6�N[Q,qL�5��`��a���mA�p#U�yȨ����2|����_�q��"Pe���QO��� e�S��?�T�9NB�~���D�#U�0*DF�@$�1VF��ӽ3iD.na�Ł��V����^_d�v3R����\b�I�ô6A��)��N �VN�3G��u����w��ϸRF��.W��b��%��i�%�_�G��(~���XY����Z?Wmr��ni�В9v�r���lI�ä���:�&\���h�se���<��"S-q�_���V�In���g�s�)�/�Qp�g�-|��u��ۧ{]x�n�l���!��v�YL�Tڕ*�rc�?�+����U`r׹}؇o���b!P:��s_r>�2�lE�����#��id6+�Y\Ź#��
S>G�$���{�ݽ6�Pg�t��ǝ3|'5>iȬ�CֱVk-h��8(�>Ҿg����~�E�Ҝ�g�δ����o�P��;��J;��CO�|R�� eg[��s��b}�1��Yeз��:���q���W-زZ�i}]�೻���P��=N��8���:��u��A=������$�n��6!�a��s���Ŭ�|aq�c��=]D��)����>D���ih�!�+��ܹf"�5��X�S�ٌ%RMt\t�,''߂_�Ӓ�Z��tݑ�MN١|��s������D�Wr�m$H酵�6�ډ�$��5ߪ�wt,j����02�޿|p9D�
7]b��j��h�7w��p�#�(��'��pc�b���;��W�Î}B;����`R����^|��ċɢ����o����$��M�)��B��R��+!����D3�=Ѐ�h.F�j#w���9��k�^>U���5>��U�%Ex�tR�M:AeT�+S/(��0Zl o�)jM��F��d���h^��z"���CZ��)��bfY�G�8�~���U�t�]�/Z�V�:jl�P���lV�)o�2ݲ��Ug���-j���b�l�/��Y���m��oT��2NK/:����Ѧ�焷�qyU/Y�Y0TD�K��~�z�F�J�2� ���g*���R���DG�F�W\��8$p��T�_�������,e��C���n;i�K!�K�cf��UY���:.T������w)�4�d�Ę"�P��B�XYLȔ.WH@���J�@�|ݻ �vI�Q�;w0�M��e�9.+1��B%�vR�#�Y;\��M�ޢn-iAi�q&E�OU���	{7�&��yCE��TQ�D�>���tνe��7�b��>�c���)7P�!��v�h'�1�7���f��K�.�!�8Z�)��7�|j� �c�vIY������)��/@g��Ţbq$��U����OUz'o����CmY���%��O���]c|�F����`�f��K8���v"Q
��Y�%Gx�؀+�'��s�ֵ��z�g/��u�9|�L�2��)�����ԇI�����t�~�͉pa���E�3xR�J��D�95�̱����0�,�8̜'G���Y;��b.��ɻ���<�;x'�ܨ*�e��k��%�2p:<~�x2U��eL�'O<G��Q�f�L����,�;<���,&�2��y�^��΃����7��x5��A�!C� ^N��f���KC2���+=�ٮ�C��m[��=x�2��ޝ"�l�DQ�}��u�v�������P�r~)P�~�ّ?�\��i���HX��i��"���xYɃ�i�e�X�ڪG�$���[ͳv�P��b����ĝ��''����UAi#2�F�[�8��IWG����7!Π�X�ۧ�:n(Z]�cu��;�WitO�Ι�p 	I��Tc�?MXG:U��)�?�Z�K�9���	 �f���;~�W�+�M�c�#�4��x�ͳ�)�@�+>�\,u�Zu��72���a�^DZ�+�?-�$���������|ǉJ��圡c���ٌɗH��^�'�6��Z�Ӌ�.JB�B�YSO�s��M��K�����W=,|!��+����C�a�PtZ��aV��[k���GOs�oX��\��2%�V�C�6��"I7iz��������<?�+���"Do�]��J�����	�����fv���bτ��4l��S��m�̼7I(6F�K��ce�G,s6[��nF��h*����^�<ujW�]ug���n������Q/X��mx	���Ȏ+)�Kn .���%���tP����S"g���}U���MS����mZ�"�.a/x���VL܅��z9��.���d#����O/C�3��w*b�{\d���o�@�J�]��R��o�*M0�s��۷|]��p]�s`}����$rd����R��Ω(�e�+�]5S$�)3dD!Q�0ޑ�H<Pc:�Ј���8�vQ�7C�%ѻ���~5�"���^~�����q��>���ϔq?����
����9֬�(������{д�}B�X���ƻ���^�{��0����L�$�OT;%���TN�a��C��|�z�\�?lħt<���4|�������?���s 8�h�c�]��	2RoS��o��T��q�L�����o3J@�=�)��0χ ��U�u�5h�!�tr���!
�&���)]e$Pq���7�Xl@y7S�Nv��vB,�łe�.���QW,ӛ�}2hb�H��Z���Ty�CQ6����c�̸�Ưw�p#��l����Vz�/YvNϳ*PK��8Fg1"���qͤX�9%�b@1�����k�]�EHvP�&{q��.�&�D��L�����m_7&��k4y�2�DA��@��+kP����%�	~İ|&�*���&k��`�;?�?��M���w��v3@�v}h��~�`GRRܛq2��@�g1U��qN�.^�^����:�ȍ�B(u�[N������n�-�&w/R��ܦ/�g�ǵ�9�Ԏ�d���p���Q�c���2��� �xeT�nzM#���U��6�rF�����!�L�Z��k>	w�#�Z�QI8�T"����*l�s���I+�bЊ���iu���=�ެ� ��������"�'/aݐM^�{;�~�p���i,� �*I��7�|n�fN��>1��[�]�ܴĺ�?V7��+)gQӫ�����L��̗{ӣ�����]���0� / ]=al󫡎�R��H}/c��2����/�P���<��|i�@�5=��Q�`�o���j:כ?p��T��}���~��m*"��F[�����K�M�q~Lnc^��U��ͨui�|^�8ܺ*�
1�)����P;.xsoс�6��[��{�zY�I�6��b gf3����|@�d'0WA��A`��� יڢ.{�^"�}��lЗ��'$� �]��K1d�ϼ����=�nh�?���X�N��~'��j���)BI��Fd�ۢ�w�¦�;�8��U�f�ߦa�6���G�������G7&����4#�(� ��HpQ[�'�Q��Q��Y���2@�.�Cft�`�tt|qo�}�Ź�n���3��1�{PBZ�@�ǔ�v5��	���x�86e�Ƹ��M�CN�����������(��Ԡ��EKi��8��*b�����B�:Q��ӡϚ<Fm��5Iߚ�g|>�o��,�lL-�E�tg��be9#�M��� �2o&�f]xlF�W[����)�ω�f��#���B+�i�]+ݯUZDVV���@��dm���􁉶	�Ī=�u�}���?s_Weې�T�U8W��j�&�Y���n��u�4{3�SCn,S5��i��:�װ�	 �rr�jw�?��s�D�1�1:�#��4��TVd"Y)��`�a�����Ɋ�Ќ�#?�m��[��4l���R��훆5[��"��0e�9��7�}l��W�����.V�7�_<>�~��S�����vv��\g]�~�r�,Ϳ��# j�3	�(2�2���l|ھ|�)=��舴ܘ�ڜTȅ��~!r���,�}�"ƚ��<�P�h�Ȧ��·����f)�b�,.��p��`�+Q��Hd��?C��`�%c����k��jʣAQ U��̱w5�a�������F=���� �4�5�N���t�N(�Ģ�-� �Ǝ �>�u�z]�$�9�F��	[�Kr���aXJM�	�8�%&C�����R���1�ȓ$���>�n�H{����ȍ���௅���r�����a�����}RY�6o~���;�o�_��4�|���{�����O�zݧ� J���.WFT�`(\������)s8�N����O���v���j�4�v�׍*��7�J7(���$B�m�s�H���5M2F�v��FgS��*L���U�SJ2��(C�>qҞ���KT�`<RX#��,���HL.��c��928����t�� �si5KZ�v�eӟN�� ����P�p�& ��u���6�SŕS4��qqp�m^�������EGycV�leՍ�[��t�4��62����\Q���*�;�u���)�|t�7��=������\F,���5o��c7?�zP!W/~7�{�ʴ�)�ڹ�)5�qLh�D�9E�[�ia�v�o����O���8���B/b��b'|�`�I���Ձ|[`ǋu�	���Uo��S�����u�&�1<�9���Z5e�M^���#��o��*���S(���p:�+� ��@ܜ���9���Jd��Cmk�С���) T���`r&�</b�.>-$��F���E9�4�<��dЋC�ٵ�H[�?;l�A�T�����ѐ�V���Յ��z1<�ୠZf�׆1���Z�����,$EB~��w?/=�]�b���r�K%��l���(�~�/����SƑ���v�Q56z�D��Ab��'�u80���Dڤ�� �w��]��]�[m{IV<�|�PiV�K��^�[f�&?�m#�F�U��no:���ئy"F�$���-�9�Dv>�=�Iyp��U�@����,��))�:c�K�M.��aOJ�p��1�c�J߲��x�p?�y�{2h�-;���X�Qo��!P��5#ʷ
/@��h���b����!�(����3K�̴�(@;w�n�y�B��l[q�柄�#Lh�d��ZZ[��c:bI��jY���\
L#e,c��(0M�{H��I;���W��~�8�,�GA{e��0����4�:�ݿ�J9���KJΩ_1�=|��L#��E��.@iѓ'�+&�!v1*6�I�D��+fzc���eb#Ȱ�2��H�b�͂�A�w�A�}(GU�u�!I�pyYs�
ʞ��ň�q2�O�塆��AI�h��d"�>�ϡg�W<�:dO� ˣʸ(��w2\���i�{�k��>��E�2�Η���a�^�]�l�쟣�l�%�]��k(0�$��ia�\���%0Yo���&	Y�ɣ�RL��JN�	��c�l9�?ך��Â-l�a5�B��j>p�]�I��6,�-�\P8B�/)�#JIE�-*K���N�?�㷏>�H����k}z������d�R��5�&�2���R\Qq�FP�o=^U�����"G�!�pkJܙ8te⹳�h�{��*��2�ѝ���7��"�5O���%�#�!���y4�)�8(N��W��f���G��4��ǰ�gٷO�i�i���W�M�vY����{��/Y>��:T|xw���l	Һ���k�����S��������2҉a� �noArtL7�V
�O��jȜ|�2�½�U���@�ba��1J�㳫֗�����L�w����W�}����T{�����1����JM.>��[���(%tu��</!A{�&�Od� LL���Eyŏ�m�����	]�xc��2+<dF�X��!,ag� GM������/O{�,��&b��H͖4ɋK�>-�W)ƀ�ӡt?NR��<:o������Vғ�:G�ZֆqGK,�A��%�ON~�mv�y��s��^���m��A���hlV�1 /�$6ڝz>)/�z�����m��}��i��GV��υ�b`?Q6VY(柅YW�!����5�ĕi-��n���B%v��=���+<V�gJK)r~�׵����2�t���\T�#̸��Oŋ�ю w�=P��K~���g�b�V�!���9�� ��c�����aq��C�x.SÇԂ�_�>�8U��$��L�k�~�W�T #��r4T|m֗��H$'8�)���!_������-6?U7�B�$����*uZ=0�A4*&˞T���t ���N��-�Gs�MKc��e��vnk;&��F�<�J	�@/ʌ�t��H;W��C�|�[����g}"�N�R8'z��^�E2��҄���1]<��/a�'t�pI�]���wkU��q:G�P/r��3��b����9�˖O��J�rc� ��J�� @&���W����Puk�X1����X�����_:d1���bI!��MV_���%@�MB#%K�-i9�������߂E���w.�gX�Ȳ1y�릖f{��Ovx���o�ñ��ߎ�.��a��I��������c}hr-xb	M�̽�n�m�f�Htq�j� 1���v6i��":ڑ�-�dh�'*?�h�\�Y\e�A:J�V:�Y C����%}'F@����C�|�|�S��w"Ѧj�"�ӎ}���3�����0<��\�`�R(����,|���/ȅ�ӡ)�NF�;�4(8MBj���P�asH=�#�q/�zQj(�u��N��<㓷`�>�L����;Aqm���`�7 �n?.r@���T�ۓ���%h�e�'�x��>$�;.=����|_pV�UlBâ�� �6ITv�w��B�9�k�Zif�~f,{�ta�6O��bF�H���P��6�� ����Gmv���KD�1$X�1n��$�^�$իSp�K�Z�KbI�h!x���H)�Eu�'�W�%�����#�@�c��n(��C�V�T����P�>�M��U}��7���?W�_m�X���R
�:��imk��QM=+�D�i���g��]h�l��iJ�"g �+mr�4�=>~&g�[�2V��j�n*�* ,gIV�~��*d��[�:���-	i�Uv[ۅ29E�\�ó�ek��L����'Jx��r�M�����ܱV�z��~A�/���Fͪ?�4u�-ˆ�i�8���wslˢ� ���|�����b���X��G���y.͡;@`2�}����8���%�jz�����;��/��ᯒ�K�SR���ވ���~QT����Rx��z[�l���+wV�k��9��Ѕ1�J��|��TSU��S����T@��V�����|Iz�z8��#��bDGf��C(1�JQRy��B��?��]����L����!emK42�h�;��������}5��u�ۂ-Nat��B�D�"@o�/�*C�:��*m�L;&���f�G����JQ�j��ha;��?|UWT�M���e�l{]�V�w}�TL3�/(�j(f,d���5k禔>��OBX��cԧ�!vl�%)쯏�ˈu��z����P}tB�g�[|=�_�A�I��;�o
�`�oc^����aM���7$cl���v�����`��g��ϳc$q+���k��^�*�B��
ƽH{=Y��j$aj�����kQM����X��N�>���}��>E �*N��y!0g�>r�+]��so,HR�}�Z�؋�q�� ������{kZ�D�֥[]5XEK�xe�[����P�5�y
fa�-�A�J������Ek��]!�����[+8`�0ܸPg�Q�~�0۠�ַ��=��h�h��2�i�_�˟1��S��#�u�����uZ��C����y���V���� b4;�-p��n�3�X�+�Tw�ֳMv`�V"Y3U]��>$������k��AH8����|G�� ��������|+� ����҉��@�,|��~��3�2�LNd3�ë���9����}��5���XN:�_*oӺ��v���臖D"W��7^T9�	� �J��F�uf�����]�fZ��b��������xk�F#8
��z�J'�L�>��9K�� �z��a����c)�!a֟�Pa�H�
"S��[�}6%NX�(�Q/�;t�ܗg��%m�f�k=�μr%X"^(Zޮ�1�Z�1D�����
�~�~Ln}�P�ssrf}{(�u��#�Q��fZִ%�$Lf��e�ez'�Dۨ}�E����{��n��.�K�dWui��]�,JiR(�$sZ�#=�U�2�v��"ǧ�д>:\J�~�iHo�A������N�Ls��
n�����UZ������%��aջN�y:��YxlV���:�lOA����mЖ��J�%�� +2���m�`�g��iD)�Ը6��KL{�:���:���Z���we��2oN�ZΖF�։UÞ��>�~$Ҍϒk���=���W�X����ᇨF�>��0�ȝ"�мh/*$%{��ϖ��"��V���(>�ڀ�k7��e%��b 7\	r���� �s��@PW��r~��RZ_��T!�4L�;��!k#"^�R��ީ>�X�I�<v���
��pO�����'����)P&R�J�䄵δ)��Sbk�%�Z!k ��zÙ�웿��.�X�i�6���ύ7��f&��8��¡*��òX�y@�F�_m�T"m1�e_�	��O �G�����;�2-k�xc2�W��/yt;���)S���2�����v���4V��7��趩7B'�m;�Bl�s�,<���O�������=nN� iW�ބҐ(ʕ�T#�4Rk'���2�>�58C�&���Ď�J1�<ԼN��=�㌇���i
��5��ʎGx:X9̪{�
�]2: �0ہ�%,����v���!�IZH�*u�G��6���L��U&��8�ߚhf����,�h=1�g�iҟ�^����`��6�O��w�.ꭶ� W,xڷS�z�4@|�xxg	y�ս#0	�;m�Y}�9�D��X�i��^�A�+��S����*p0�ٿ";����vJ�nu���To�K�Ƥ�i��p>���^S�I��
�� �T���Sذ�iLH�:�-��%��.�z$�>���+�zzD��yx�n��GY�Ui͚.RJ}/ �U�tJ�-��"�R6 ��ޚ�R�p�EC-�F�.��/N�
��R-�]��*���Hv�Q;H��A�IZ|w�B�f�:L���4xK^S�=:�#J�i�#�����r"��_�8����+nx�!u[Fm�aQ��@b|X��\��U@G�!_C�,<�"��d*;�	���-��g��尙�}�RK)�g�MSQ�IXa�c��\�6;�gʺ�W_�(7 ���{<(�ߗ�����8�¾�OĜ�5ѐ]����b�$=�2�N͂���{����<"�	aA*�IXz�*_`�R6��Aắ�����Ր,��\q�Y,�;��[�������~�V��Ș���i�7�A�鎱y���yj0����"�4�x�`�ּ+���e���9d�G+a`��0S �iP�3w��E5��P��0f�c(T�a��번��K-��d��S�{�?��R�bA�ݟ�b'�����҉\�Jq�Y9�f�E�˔<� �]�)ҧS�K����h$>��ېbv[G������bp�YE��Q��#U������6���S�\�[��q��D�|����#z(��~�fX ,�Ki�8��`#A���uo���������4��X�w��B�@� ��n�==�a�[^�ʠ`i�&<��BW3a�Q�ϲG
�.�y�ᎆ)�|ߦw�zM��2Dk���I䋀H� X�wl1��Z8y��]�W�JE!2��G&����(	�D�Ԙ��]��X�R��~8veK-(˚?���&�� �t"$T���By�v�K߹)���Y5hA�$�e�L��'}.�B-�U�7�o'ᄻ��@B/�6���{��+����m�����	jzw�YsPH㕘!ߙ�!����N�{�e�\�#l�c뵏Cs`������7YY�/<z��+`�M��iC�����QV�3ݵ��C�t=�:��g�H9�rz��#G	~��'�	{��~�S��B  [I+����i��Hm�j�xN��۱�xt��_��yܰ!8����[WF�Z�9��J�� v�w?>-α�
���úXZS��o׺����������C�'P\�j��<����d~j���Zp~�^�+��9~�i� �_�q��b��(��TѧBc�\�	[�B���P��5�0���$��mh*J]��U�s�(#�_��Z�F[���>�P?E֞��_#F�q�C����VA`�;�DhD�HRz��γ#ڒ�����������IE��oT�/��imIQR�X����J�����H1l-r�d������<юMT;�!��dr��)�,v�j�R7T��2�:�AQ��L	� �g��_
L_���������~� x�i�/��c�D~��t&ګC"oۛݍhя�����4O��%Q�@A+G�ܥ���ٕ�uN���@l+��Y)Z\l�{�ا�&7��1m����ʽ���[#Ip��]K�S:�]���8��3�{"q�P����*��5{���P6Y�'�+�y�z �!��A��y���F��n�6�����X^
a�I�������>�ui��r��� ��uxD�v��lx��bO�{NpN7��k�O.�~I6 K���ip6[�J�h�m�8�]c��Ʋ˅�#�M�-�Q�"��%n��0�ϥ3Ӓdn=�]}�2'��� a��R�"�z��u�ǎ��	>�Z���Kp{^�餺�����f���E�F��˝mQ:�Xt�av }������,����z����� |���Ӹ|S�Ӫ���(Z�K���.I�6E��Y������\]<!;�\�
���e�LL���[(dV���Ⅸv��{�U�n�x��~la9��]���SR*�Q���?�W�>�_�6�0�\�"� S��Jӵ��?��	��M*8L�0�ud(sQ���3��V:�P%���-M��$��Al �����Tu���)M NW�g|���P���2+�G�y�^:�����n��Bv�R��>*���@�(�f�װ�����+˦�f��x���K9�Í4�3�YD�L����a��\���k�â I���t)O��������i����"�>Dp�)$�C���mY���������rc`�^f�Ct����n??�'z�}2u*F���q����{��L�_a>�Ud�5)�V�L��|�J&/�P@��|���{�̈́���0��I���`����s��-�3�7���y�R�U:��iÚ2���J��L޽��=��9��UOn@��^�tf~NA�U�J�:{�̹Vy��������$
6����	gVD���������;�Dm�vCU�����[��Rj�͐�NF��=�t�p\
�ٱ��xJ@�������C��b���>{b�H ���>v�e�W���i�3O7�sϟx�ׂǸ�7��̇G���QE>���yP3�0\'����У���0��$���V�E�����H�nG_6�=�)X���n̼\`�����?����2���������ΜS������q(D�dL�uY3Ã�tgx���L]do JFw��`)0�)o׾���Eٽ���o~a��­c+�3�.;�"R��?����O���E����&��X�_V�C���-}�8��b�`CsK���h�<��;-�azrjհ���v)*4�[g�[�Q�^��¦��6�H?�bQҳ�] �tt�	g�>/@�3E���L��H���\�&q��2�.���a1��������Uc~э��T�u�E���(�p1 ;�y;QY�4�z�#a�-4�X�B��*2��zC����ʨ���!t0҃+�����< ��C��3�+l�C�f�*}��=��$�a�=�(��z.6n�	P46A[,�cڎqx�uL�33��z��c
���o@�?�`����3�|h�x1"Q����o�� ~�	������A�
�Qd���k�Y�*W�j=e��3���bE8x>-b�驾w�Ϩs��\�$�,|u�)���N<Ӫ=O�`ػ���(��Z~b/5rw����)��tU�AL��?Dlo�p�k^8�,�D�,z���D.ͯ��C��W���}�NdH�ևS{	��t>�_m�h'��ՠ�����@��35Ô����:�h<��";UV���J���>싗����&�R-_��B-I>إ��?�C}��W��>)P@�YH���z�иK��UAI��r�jx	���x�Vc��p9���+��� ���M�V �]��	]R�)
�1�k#z����ז��9�Q�lט�����Ve-!T	����_d���]\�2��k��T�!��9��v�Bo�u���p{B��[���7(�Pk����26�n�������U)1|��pM�����\C�����}����.��	��$��י\��j��u�"V��w�L_��6�l���lL����o�Wſ�[��S+9+B�1��ݹ�����yA ��bvE̷�j��D�
r�{K��q��뾘c����ȋi�i�Rz���� �=+�9,{�/ ��Q� ���oi�!�`ܕj�MIZY��J����̴Zd\�W�Q��2%����
G4`U�8z<�LjM����6��1��s����rXZv�B�+h�M>�G�����D���2	Á�/O|�dP�v^:�JY)Vl�'�u˰h٫�;kgb�?^���RζD���5�Z�)�n��d�6O�PN]Q�r.�g(���s����j�E������|��;=~[���7Z_��uz���P�3�6AӖ:��&q�\�#I�lm
%d$�g�ށ���T����o�f��y�3��.����j]	W�dʏ_J񿆛b�r�>������8��IpF�1��Gj��;��!�
zSʦ�G���'��fI�5a��=�5 �Z�Z�뉋�4�,��I&a�Ek�>��=d�؇��+IJvH\�6��LG������ǔ�������Ѝ���'ç,ؗ7v��`�$k�e�_=2�1t����]'�z��&գ�u@>�Z.p�|*�'������#�aQ׍�Ю{�}J ����w�Ggb���o���y.Li��"@U'�\1�tF�gp���o��f,24��RI�^ �^2QO2��li��i�'��&����Ȉ)�2Z\�u>g���J�˭X�9[��f�ߨ��_�>�i��VL�	Ц�D`�iɨ�Q�@ݪw�1���	{�Jӛ�b�躴6a�1����C��7"�7
�mR]k�"9���B��h��@ü��-��K�N��ҫ��z�F��K�V�wg�gK��V�,�����Ɯ3�'t5���h.��-�$?�]����$,���G����fO��(������&+�A�+ai`9� ��^��&_�WTϏqe����t��E��T�����ړ;%F�	n�Z�h�
��9���Or��1�Y#�?�`vf�_���r���7_�Y>�㴭���zj>~�0��C���W[��N���̟�H�ݒp�(n�Gh@�s�/�\�L���wF>��`w�y�y�>�e�E�q�D2�o��'�%�b�|/�'��_C$�)�����w��A��W�K��CJk1	=i.��W����v;�=I�����)BM��Ͽ���<�54�����]u�m ��$J��u�� �$<�^[�b/!�:���.{������K�(��|�`�M���,8�����&Yz����_���{��:*z��=�KU�Z�O@R9��ѹ�r����9[�Q-��=��MJ��q��SZ��nX�ݦp�-,_`�L����T;��B�ݟS��X�6���F!uè06�]���
�!!�t!zגݰA�"�Z5��s6�عϦ�F\���X(Ɵ�iHg�ˉGCyr��9/Zpg"R%��RA�bt�~?6�̻?w���Dm���`��Mq�g0.�,� ��	��=����~�r�s�� ����� ��B|��g)J	�ZM]#^'BR\��q�����Ս�̢���3��Y�ܠ���� y@��3��=j��n{�WY����:�4���ཅ��w{�<
�+���\�iE��G�ub`3���`��R��ɟE�&�=�uب�.Ns[7|mu����T�)If��$��4��m(p��(�xa�R������?w1=A�9L_�ꈌ�O8��)�lJ�	�p�9�F@�L��Y��jZ�Z��*��Ƭj`�����vA�&O� ��c@���4�1��$]�P�f1���C���*���PrzM��}Е. =������*[YYZ��HD}�����%��0��S�G���_XT��9�0�v����f�n��?d�9)���i� �8�C�����G���ǔ{�ۜ��y��~�A��Y>��+}yw���r&�Pn8|��^�cj�l�ꈤ�?,�G�$t��@5'yY����fF$��d�Β`�S�X�5�:���ك��*��!�P��^��j�Ä���rfZ`��B�d��"1oV<��y�\�=�Ёƌh%5�Y�S>��5�s��V���+�yG,�|H}�s�(RT����q�y��1=|AE(ל5U�3�"k�e��p�1HN|0F� �e��,�l�em���C�K��QEZ���ea�c�r��g�\�ع�ʂ�O��,���K�(�n/k�9nTzu�µ������+��+�}��XF���N�="��]k8�������_��b� ���٭6g������f+Ǣ�^��̪A�+�Fq��Wy�{��%��iNك���\����L�?�$���i9{?3�ʌj3��=���k�b����vt��˼�A�c`�S�������7�(����2��D%�������̨@8�����P���h�V��0z��Y�)j��l^��������Pv�/!�-��u��� 4@2�q�s]Dt�]Zy_@[��a������đ�a.{����0�����@>Tݜ���m�\͞�t,о<�v4���a���>Qt��;q*i�'x�Mr�[V�
,<��#���>[�M�UMRL�$p`�f�%����SiQ�@U������P�oE�'�[i��b�JR�����
O�8�Ã+ D�e�P�+��x|l��]:u�M�A8�֏Vg��ca��礹��=Ӊ���Д�@�1����M�[F�@
<-��`e�'�Y��YI_��1Wu�T��؏��l�������H�*��1��Ĺ��9ᢓ���ȱ.����	�Z��{�`^.`k�#������ H��N��Q�f�,�?T���p��cwu�����p��'�[Bs+X�̨.I��鳃���V�QPp¯V%�����}w��Ȝu}�Ov�=�bGV���Fd]5�s��|Z�\L���_&e��a�oa�..-MQ���^���6k�&���3VB��C+�G8�����+t�J�X�yZY��j�l��&$/Cތ���DB���R�A8����P�����N��S�"ET��>������<��R�NDل` KA�ğ�C�����Z�{�:E�SD'��������f���F����@��D?���U���*H�����c,X��&6���7���x��^�+|��8Hq��X(h�~P)��I
��D�Mt[�y���#�5.���{�z�x\83��<M:Yѝ���V�Ɉ�0#���߀����C �0r-���@��)�����8�.;����_�s���8Ҙ�&�/���*@q����C�N�ѧPY��&�jJ�I�,B�"wǼf��Vk蒍�0�9��=D���9��g����#8S,	"���:"k��(XZ
�Q6�c!e&wtm3	�-�wՅ9���y��ށ<+����7G��O��Ԛc���*<Ԏ�9�sSp����e�kW/��(��/��g���5h<�p��p�:���=�bNP�����wK]e}cGOTʎ����ie�����Qt>��SYh:�`�俔��ʃb#R�����6�Wdꊅ��ۻ��;}�t��1W�d�gg8s��8�H��A��wąk���~+oXw���TW��+g�S��K�6>/�!�Pd��!��
�r�hk`���������'�Z.!�)�¶�F���;��:���)F,�6�uw_��4��y�����0���*  ��YS��K�r�>Y�S�A8�*�T|?�/ӂ 1'e��|�7�����X,���@��Za�$��'��h�M���.���^!�{H`\_�~g�F��~G�z�jU��J}�#7��k�XR�,=��v�������:��hBؕ��Nzq��#NI���ҽ��$>�1��A>4p�������$)��f"��8E��-e��#
�o^J���Nb@T��P�S�_�m��7�,D����#[�KWTw	;Ō���|�?�]PP}����0�y�*�¿��+��"��\�{&Y�OC�cp�E{�I�'cWOzNStW����ȃ��>5a�p�Eǟ���>5��}��f!�{�R�mZi�p6=��8�!�AlD��^R�������:���rl�C|��@�M���/{�R�Z�5��,�P�I>0�OZ|��"84�	A.��/�{ړ���s���S՝��#�;q/i�ȳr1�,I�M-p&޴���Kp*���ݳV���K�g!0�BX����UZ$��&��!�0�H^�����������㣛����MQ��"OO�7ءR��0f�UE�D&�8��K
gez�;^I�h�/ц���J���r��2j-�wP��	�<O؛��߸���:��&�����Հ9o���$J�}\�:�	1���Э��c tQ�Q|��4�[�v�L�k���Y�=6�r��}��q�t�� -e��2�&w$'��HkCm8'̣W	�� �bU+5TlDx�^��S
U*G}"B�Q"G�
s%!q�´��[�I��M�:�����׵�O���L�A�xP�IꨉtV>�f��QFf��Mo�#(6D\�r��z_u6�$Uy��髧�fV"	m�S�uC�Tubc,z�)�T�5��%�{Va��L������O�ϗ�;'Z�D��e�O��ݛ�I���Tl�̸i��F[8�k=A�����Cټ��W�`��	��P��3W s�yr�4�=yW�%O(�c���$�g#E�(m�n��㶱V�=� :��nx��A�t[&j����E&�X���<��`�q�#��:>JC�������p_ x�����}���U�a9���KS?�%�f��vҾꎟ�p�R�-��;�D��2fh6�G���Z��
�ۈQC.�������k���h�^1�>9^��n(M\K�1�<�%�K�[��-B���?�\�W�3eN�3�+m�[����=���|��)~NhԹ����N����]�4x�4}�� �3)z�;�5�E(~�'"g�{͊�jG��5��$�7�P�j�:c���lN�EٛV�;7DcA�ա{kѱ�}0a��<! '���.�"X��.�K^mC(i��S�2T��?�N����#"�^ŧ�u�q���U�q�j�$�/Y���+��TC��SLHj������M�f��ݝz�'sV¦ʔ3��πZõ�u^R�>"A��!'�o��y��Tn)�0����;�bG=��͛�;c-H��Vw��a������3��sjb �7�$��מV��
�]�q�������F�D�Č�w�( Z����0�����P�8��nwބN�6e՘.q!-���$���P�4���S���]�e���C:nf�)4��	��N\��?ޞ~��bQ��ox7����a��
����m��@�T,�W2t���ڭ�ԏ�YV�^�d�W�xژn|a�WP(�<�C���8��f�����&FƙeD�Z1�P�^������sw�:��X�%[:��y��>Ѣ�� qW-��m2(W N���/'��������;G5>���kↀ~���U�Sw�@��=r&\��zߪP�Z��L�PY����\ɚU�v`W��A���]���lj�XX�Ռn�H�Ow��(��R��_�p�q�0�<�>��M�d�W�@=U<4�3��ZC��T�n9\T�
��-v,Mo������8G��1_�� )��B`TE������(vh����kWlr�=uq��40y�~c1���J�u�a>�����o��� �b;0 u_��s��,��~"Sbk@V�`>7�<��t�;M���e����&,P*�s���^KQ(��P�C��#�1�cf,�&P��l������F>���F�xJ��y}��L�?>�������<t
u����Խ�ep�Y
���Ř��:7�4�ܠ�������*�
��N�t�W��JV�C6C�W)ny��7�TH���ᘸM"�tr�u��=����e��A��	ҿO2!A`���B�E_o���t�<x��V$p�?�~N�/�������`ӈ�k�7��5�.vJ����-��@^ͺ�>�L��uQ��ң$PWd��q'� �0Bd��"�׊;
3P+��4β{�h˻ݾ**���J�ĝ`g��N��f��;�a_+��/�d�#���9�AD����_wW%�Aq]�����-�Y��F�T�[��\�qs�hx(܃�q�A3~VH`����z�Ŝڼ��� ���'���h�^T�A�-�A@tmPE��I{צ���`GOL�_Č��N_�w?mt��>�c�u���{�6��߉3JO�]4�Q�(}%_(�I��Z��Z᫝:��dGc���<c��nҽ�v�;W��VPf4�X��"YB$ʳΌN��{A�*����u�El�"A�I��@��r�c��%���U���`�w��>l��̈́��̆��_W�1�iG�Y#�p
�}iWf�#���t�T�(��j&m.T�:� �
��nh�P���p�e͡�P��Z�l�ߤ5�����q[jW�����Ѕ�q�<w���-xp���b��_�^�bL?�+B�<�[
���c)lcF�]���m���OC��oٌ��ť����l��3��ݚ@`�%��B�5aV�R��@�* �'�W�ב�0�B�n-2�r�{!����N8u���r@�P���!.]�W��0�H�S��T>��va&��We����H��2]��3�mFY����M*����YK-��m�ǿ��_V͓�Չ���G�̪p5�0��A*��(�+�:|8�&Y�2��u��.G���r����My��cU�d��]e��<��-r&�g�Q�g����;7�ۼ��_'2��N����r�,�5��� �x���(�Co=(��\F,F^������z�֋`�(��^�R���<��)(LA&�
�PDO�f�t_8LO:���e��X �|�ep�|P�'���Y���E_���e�V�@�����ia.��56B3Z;�t��Ӻ$IS���e���*[�劒�b c���»��I%�Z�O�7��Ү��Ƿ-��9��}y��O>	�=t�!%[�@5&�Ӽ�n'����G�`H3�&	�9��^����&V��,`�s˲�:��h($�;���;n����<��h���~����K���?�P��a}�0��Aӈ�(9 *?1`��J��͕L9{*�{ɟ�=����0e�j������Z�(��ߦ@�P�Gse*eR�P�?c���􉪤dX9�����aB-����&ى�%�kw�uq ������x$��e�l
䶒�Z@x�����hMnfmd�(�w� �$�z�L���x�,�-���؅'�]�1*�d�Rƌ~EB��O��Q�^L�j�(��h'�����d��o8I"v�M�X�Ż� �E���=�c���w{��r�Ҕ*0Zd��:�V�99N7����=��C�i�5?)�ek�5��g�d<C0{ũ����S�j�hH��t���4_SBc�I��ǐp?�;�Զ���J�7�ug���B�O�ɠ��?��ѸVɫ:����.΀���(sڇ�h%P�����r��=R6B�檩�M��Yj��C�-�^y��%K;�ÏXM2����8Y&�#�g<��K�����|/��21����������;!�4h_��B�^�R,��D[�t�^n�S	��O�|�?�,� ��:�������0�5�5�X���w=�۴�WG�����w N
�e�U�%]�u��V#j=�/�֛��g+��8�Ԉd�=�W���wp�q�a�1 `�x��J1�����H�K@�j'3��a�Be-��W����0e�t��Wԃ2�����!$�a���b˲D}���sP�r����������ysK�b����=Z��y�U-�=�M��4{�Ȅ�F�i�Gqha��խ�&dA��z:��t�'�߰Ĕ��i@�n��4]��us��I�q���	�k�jO~X A�b澢`��h��m��4�݅�T�'B:��}����'k� �0@XUm4�7�������}B���x~Q�{f<�,pi�Ͻ�f=gJ�����[X$�yݜ׿�Oq+-�g
p��-)�Z�7K���1,�0��\�uo��K�>o8��K��c�w*L��{;rP@�I|��	��R}��b*���r[�:%7���s+�]�X��|-�v���St�}(�}��e{���(��md3$F0���7'���)��眧�;� ��cM�zH���Tը�lH��A@ǁ��q�ٙb�pT+C�b��;lF�ga�Q��Lw��I�o���!&�mOG�[e/X�6��0M������ì��&@��Q��/&��]�!�LHon��Ө��S|��<S��/w��ns=�4P�:�Z�zc�z;��gi�+���G�y��LK�)U�+��\�3���>7���=W.d/߹�O�~k�D�c���cD^dὸ�
�v����:A��-��ۖ�䋯2��W�N�k����q?���^��zъ���J���P�
C�U`�����v
�_3*��N#�k�@|��m��\���V��n��8�*�Ƚ�����dƾ��
�3�pA/�^(�������o�/na�d��h݀�z����5ъ�%��a��'���P�>�ߦ��'$�!j���hj��8��r������0{��eMZL��p�|�q��~3*ߚ�����j/L�G�]�%��I�P�SY5ז�nxT2iz�X��6��7�Ԓ����$�ɼ7�v� ç[��� �
�ۇ|�`K�?q�~�S�:R
�y/���d�O��}T`�Wa�Y���
g������c��~����0��(�z�s��~8��y������zcE'���w� "*��?�����@OV�?/f���5j?]`O�:��9�rnPr�^r/�H���m�e�ibGa�맠(����&��A�S~�!`f�х�z�]�bM�"p�P�.��I�SzFy�7�����;�H�r*זu�H��Z�㰬��f�YrJ_}���ݦ"y[Uq-�2�	J�2w�S��i�%����S)�-OF @����my4��;����M���b����d��ދ#�S����:i.W�t��:���ixV�K��K6�is���Ġ��EW��yXu��q�S�gL����BD��B����ό9����h�շLRt�u�NNa��qfvz���9Mt�� �X�K8�(�@x����?������^��Ɂ��~{dz'J:�s�ė4(�LKy���A�V����q{;�V��X�B���k�HW�A�Ez&�JM���-T��1M�y�I�$Z��PV��\!�hC�U������dʒc��&��GQ.
g��C*�*�L�����K�����v�2��=X^n�;	�=���T����qc��>	R-�Xc�Z:D���Dׁ�N6�*�J2�i��w�"��'=g2�o�À�	k~��_׎П�H�6���H����thl�>��q� �����ݶ����ؤ����N/��6�d<oeznz��D�X�[�E�<��T3�:l}��6�M�yCz�w�F�!ge�l�>�ł��1�i^���|�ΫUw.�E6�2��߈@o�x�?��/���{VgI����v��@���r��*�IV0B�+��ʗ=z�d�8�S
�;��+Ta�zCN�n:��/�5���<�b���QP�;E�>;�����GZOst�f���}�"(^F���`��y
L����f6r?��jw_��
+v5s]� W�ڣ��ĭ���B��>h ex}
}4��5����s�|��h&!0���I[��l<�<2�����H"Ց5�Hk=,iÉfvo%��{e3\Z���h�	�;8+��q�3��F�h�r������ϑ��h�ք�O��<\�'�¿`A(D�mi�2�7O�K�	�"po���!���Yd�( c��EYS���2�gIm��x4��k�"���Vaip�2�����*}�\M���Nk׿=�&'�m�B޼^�D��fÄ}��^}�l:2�i���Z�^-:F��D�%���li%N,���h�%�݃�m
�.W�f9���ֵ�.m
���bw�0g�d���-4�?K�ʉ���y��{���ŻN�u�
/�;����ɼm�Ԏ6�i�
�U�N��l�k:�i�v0}��쨉��0��v�W�N)�ǅQ��t�xm��H��Q���z#z"�<?Ԋ1���k�����'���6heF��S<����U�2��7��t8�D�O�T�Tbӂ�q�G��߫X߁�1#r�>����쑦D��%s�4��*�;�J�hl�@�("��=iB�����*��B�(Lk&��G�.PQf^&�7ĜR�"���������l*�8W�*�4IM���|}�M�r�����3��Q;�G���L<�n�b�.�ś�v"s,��+�q��(ψ�U��O��p��22Q����8�C�F�!��u)t:zy�l�)}��l��:K
��moĉ���5��?��Ȉ�e��|���r+���,���+��d؝�k~�� T�E�닎s��m�V�� ��� >^o���J�:zdY5C��?vU{?�ud�t^Y)���0s_�PC�� �W ���΀�m��]��t�����6�����EBD�oX��M﯎\z��U����ޠ�X?6�ªճH;�u�\�b�����s;�H���)�� ��[R��UW�
��@��	~�4(0h����k�5W2�}�ib�j7%�����e��7̇{�D��s����򡸨N��GH(�X&M�^�]	�ӔG��W<a)���� ��罵�����gGm|"��1�P��u5�oـ$P���拾o6=mQ�<��h����}�!���J�͆p�R]��t!Xt+H�e�b~�8�A3A�*)��8i� M-2i�l��7�*�Ũ��߹X3^�����`���x+�>�T8"�"�����U[��gB��h���ˇ�|�� �>�����%�|/\)hCS6@Q��V�	�Sg�� ��q�f, g�9d�:��A�X�����+�S�KO��h�c9ea���r >�4����J��ui�4�b>#=?����,��;����:Kw��g�BG�S�S����0g\H%s�X��e��X��_�uKּ�r��*����%5E��ƨ����)�h�f���0܄�0p�E<���S�����{�ۻ�����Y��LK4R�ke��/�C< �k�O|�A�%�&�[=���s:��$�0��M⯫��7�[0�l��&3ޛ��*��k9D�O�mZ��&���Χ�ޢ�9��tvLɀ�xvZ	�H^:����~i��ӭ�瀁m'� �:��(O��(ÅeHW�Zs4�l�����]�=Gvg���
��N��S�U�	y��&x�G�ɾ�2b>�nEۡJ8	��<5��Iv�>5��{E��y]�� @ ܂c4v�a�ν0��;�pJ�
��%$*&�xܱ�6����Q���"ө�2D�($�دuB0�%�T��_C4C�
��E*f�֗���݂qb{�̙�HL��&
�I���� rg)fu���3#���O����n)ms\ڻ����Ę6Y("�ݷ�^�>4�0��q�62Cb!���E��(%�bKU�D������R�x�8ʰ�1�#�����&*{oo���έ�	�ֽH�����a����DlM�B��3��Z<s���5�hd ��Fv�Y�V��0�������������6������$�_.��[,#�!��{zX�-�:�^+������O�ֿ�FO�K���5��*�BcI}[���"��H���n��G���6 ��۞�a���#ܯ[}C������z��8W��q[u�W��҈�&���SB�ǌ�Q�o��Fo�?��"�$C%�75�|4C�d��#C����;�ژa&5�v���0���r�ܩ
}��k�<5|�i>Ra�`��'|d��?3A�Z���7�:��i�����c���~!Z�0��Z�°-�o]�Z���]yH��d�SS#���os���<�+��^��Ua�����
�-2���p�߃[����N3���l��-q��9]v��{�7\1��QT��^9}����Q�`u��={`G�OU����6���XxgŬ|��Vbp�ߏ����51B���nÙ��k���Qش���P���\�>�`�wc���#��p3ӏ��ڹ�}ey��8��������P~7l>J����=�P�_�7:��B���5c2���vǖ���ɤ��*okLk0�e��`��·�/35��{�o���������^�Ц~6q�V�����,��?�a<�͜j�L��/[l88�.�]0�蕾��!�ấ[(#E)�$��KO�
=�0�W��_݁al�R��>.��1�<#e���n�ɑ%�<���S0���<JkI�I*­��=;���)�+Ջ~�JU�����Sm;M��H�^Tͱ���1Y|.d먷�o߉�c��8��{��<�/�޼����Zib�rK^�j���ɔM/��Ҿ�:]��c0���,�O��yg��B�����%eA�#�e��J�����+��_�
��lm�3+�j���Ix�0��8�azq,���<v�U�T���1AB��[�hiI�+}q-o�3�z���_E.���oD�\w��ǟϥ7>������_��$g���VɼF0�0�q�;�o�F��5�(��[K�f�3\@+�_ u��]��)J5����u;с���>XJ��ѡ`q'ٟ��D�0�G�E�t�`�s� ���HI���o�c��p�&u5޹Ir�L�3����o �#����H�]M����8�^Y�!LWm)��a"M�T�gӁ�+�y#5)�d���3�%$���.qt����[ك;�9J�Яl�>�W����#<l%�m2T-��O�����n�Ӑ�9[�@0\��g}38U��(�o����Y�Q�|)����Oh�25S������3\��s�W��^���o$�H$[D���������v��8�$w�ixQ?��e�(5˓��E��q�wRBs����ȳ�9&��ʁek�p�%ßD.�C�{Bg��<���z�1|xN�I|cx��d���4��u��I�m�&��૥h�D�ߒS*����z;Nv��!���V�
��07�1�%��:}f���<���뇎ʽ�O.
�6e�?�3�����.������=�U�t���j�fR�̤["6f��k� [��z�]���ޭV�2nn�^#��������F���� )��/	ۤh�K�R�#x�!t�&��B�=B=��K#N|�]R:��Eo�ke�r~F+�j���D�)��p���(m��z	Y�m�(0e�-wf�n�����tԴ����{�E[oC�]��Z.[�6��� ���+�Θ1�Y�!�)�2`~�_	�j��m`l��t�慾�VP�H�Ӓ-Y���,�L>��>����-���������mce]���bLa�n\�4����,k�';މ)��1��f��v(����_y��V�`���B�bl�*d���NQ�	M�{�D�o���O}�)#����HV8�=>	AH��"�tq|�HR��v=��4�ˎ_�5�o`gD�c����XQ��b�׊�#ځYš��13����Cc42�j��]j��IT�5$��z��쐌}�ѡR_"��	B��g	�}����Z�l/H,ά��ot�v�n����Zw��������d��I'�f��*�ȵ;��H�M�i������k�^K�Ŕ�a�s�Ӛƅ)廇a�{>��:j�n`Px�Z9��3O��
$�~S�p:��KL�A�w��5��1��Ku��h�
W;RK��@g�fx�A���m����� �,�Ց�_�#9�(	����fy���4�J��z0�=`���rԓ�q��C����R��8��4@0��!$���KTL �������m+4�K���'l#��P�")a�yY\ԓ���C���n/�/&7||`��L!"q�Cg
TR���T2��h��BE� ϻ6�ۘ��'K2ӟ��\�$2<��^���{�).���@�[�%������zs{���fniFH.{��-���M8*���K�u�,�l[�sX1I*��t@�#y"Ҭ o'f��� ��tLX��s:&̽ݮM�<�CIj�7�����T�2?Ն�,@B_u���*�5�"&��A����h�JL�;�@IB�Tp�qd��+�,�.k���oh{�Ƞo������+��7�a��h++�xV�.ޚ�v��I����+�&�x�>}HT��^Y9��m����]"PǢ��`�Q���_:C�o�֟��RC�dw*� ϝ�����A��[���&�;����Xs+�x�-���ݐ���P�fy�0 k�K5���/҃,����W�����V=B�z��10�����;�y�{^�H�E$Ӿ��
&�Y����|>�7�����h�cphEQ8i^��`p���Q�U�3`�\�m�T_��[)��V�w~�/���������>���_�����-��swY�b������6&��a��BLޮh�
v\��q3u873I�g�D��\�}��d�-Y*�mu�H/�\���o՘����(�5F-����e�q ��L����f��=daC�"�M���4HCy*�H�n�J���y������?k��cb���\��wA�`��^�ٽ�|z8K��n�x$}�|�.��Х�n�p�G~"�ͬ�^�(��$6mi	T������g���[�iC��j�q"���Cy:���g���
ɦi����E��xOQ����	��M��{\���u�ZB��|�J���� �s�w��M��B�ws��\v�<�(�o��T�����6X:�Qa���8��xBw2���E�[�,�^&�\j����w��6��ւO��-�W��>�鈲	3ƚ�Y�nL�����"�%]���n�;��� n��>�1����^(j����H�l���H�G��A,�>L6mN�:.��)^���	v0������ y����*t��(��U6V���[�5����u�x�_`�׺���e�O�;��5�7iC+�M�����7����(Gts�R����k	6/@]!���q��b=�{�Ӈ��F��-?\�^����{����ȴ�J=��)���
��,)ȿ��PyͿ\����*Y	��)�-G�ؠ���<��-��,� <[	����I,�?�|'J�M�?6Y�g��9�ɡ���MH�G6���O�)9?�1G��{E�R}s߷����|R#9�w��;���}�c�	?ܱw ���uː
����r|K6\Nt������}��>�<l>��O���@ǰ	'¹QF=��YW�O��N�*y$�P�dK��-��*yh�������@V�˽R}m	��{_�[^�0�F\�l�S�zK�j5\����bu�������Q&�C�=a򘜁Cc����%���o,���3Xv-�Zg����4ِVp�`i�Q,fW���b�d֥���^�Lyf�5*��| M�u��ܻAv���I�|a��՘�?�˪���;��s�\ƪ�1:O�\yp�:$�[��ў!̘qT�5{^�%*(�u�,N��kc�rC������|ݳ�.������ENZu���|�L�+h{�	m��ĴAɓ1@^3� �t.������.}�\<f�3k&!VW[���]�cz��R�J%������'���2����b#�g�/��64�3h��I�/,H8<4�V]%M��}ԥ��-�w�@F^Ðةly\o���0w_I6��N$�o�$�n��M��6�����v2�O'���j,
��$�C�)����/��Aܝm��lb� ������H���+����4"%���g���xBJZsv�<�(�w�>B�2��X���L��IK���<���.8~���a�Jl;����Ù���Ulq��cB��/���G�G�\EŇ�N��U�P�.+��:í�@?QU�i`c�uhV�����X���5�B�޷M�G�O@K�S�.��%z�G�=�)��ێS��5	��hn��L��/n\��!��Y��zxH��T__�fg7hCe�U��S�?fW�P���[�wRB �/�!!]����Qw�4J���^�r�z5=�^�q�pqy��x�����\HV��>��݉Kj+
W�}��eh�)=�a����#E$D�p�D���2z5���z'�m|���P������d��xc�v�JyVt>���2P�]d�d��}������	x�`��g0�	G)a�Vu򆈟����F��:�}!�M��s^a.f˻��x�F���Z��V�����r{�� *�W���N��һSj�U{Z����|w���x�/��������H9c>��?�,z���"��,��V��D��O��r���x���;�F�ou����2��.c���4 �X��~2�����7G�����yYvC[����dr֠\����y3�}�[bamg�у�ld�]��l,������7�/K5AHM2/4���c��5��r�T�׺����a�8Ryx�C>�ֲVz\�LK�?G��k��������^y��P�q��?�B"]�ؕ+�*�=�c�X5�l��-��#�]�����W7��BgJP[�� �=���L�驖��:�\�����z1P���酾R�T�;,/=������B�_u)�=�C�[�'��+�X�c��[�*�`v�"��T���a�p�����Ei)L�o郻�̡a�+�-+�%���=Gս!�/W7����T�����L�j��]��<~�~ �z�u�*�g��`���"4�\8�tϜ�:|4)W4���O���1o���� ��qE��^aɑ>��V�2i�^�X�G�0��ۏ
F�~@k~,<H��n�RU�/a�m�wt0��
�QK����ն�jgk<�ֶ�U����Ѻ<$�8����ȟ��DU�O�w��c��A��A���ʛZ�n�����ͷ�K�(�OJ%�ڧ�LX�2P���p�o���'���kzt��������k��(��;���9���p :��W�� -sǯ���||�S%�"��C������ҨĿ��{�<�P��u/�]�dq@�R��{W|N�#Ȓٺ�T\�f�a���F?�閷��[M���19�`�:]A�+�%Ӥ6��b���� ��kssu�B�\a�E�ũ�Ӛ�6���	�?�KLn�ᡘ��`�*+ -�v|*,��8����e~��[	�o���IoC�r<���>Q�;)UHLԜ���k 9�z��dE���fAH�|�jv«��
���:�*��Z��L�iP��ʸG+Ѭ�R2�ߝ5����į������~��n�n�Р�T�hK�t:.���E�D���`j�u��N'���C�$Q��!FؙbZ���q��H��V{D�t��Ի�EЁ}��#;$�6$��6A/V6����9��_e�@DfX|�m3��q O��ѣZCRK��빩���ȞH^��t����ꌭ$v��<�bƦ6�bs-��r��N��hP��;K�c�f#+��9xq�����K�iY���	����K��7���F�{*$~q7b>�O�����i
3"^�Ԋr\e�������s ��bջ���>J.<�ȨR���ð\���/;ߓ�:��qDj������3�(:c��{�>GB�s�^�\7�-[p�p��ۘ�b�J6 .N�e�L�b��187X؟����������X"D�v��&�d-6�����`��<��yP�F��eݶ��&�mc^_��e�rƏR%��
�����Z���+]1��V�-5>����AV�~R��S�О��z�أ��lp��:��V|�������*�F���`,j�1kP�&:�c�E�?E�"�]�`�1i��i�k�6n���
�$I�5n53fܣ=��yhzm3�g�dbVٵk��#Q���k��Ng���cLE�do�ɒ������aO��ո�<AY�c�c(0;��#����j8iB�/5?��ϜǘIPj΀i8q��w��$IlF=H@��Rڵ�����	�C�ײ�Sh��١�!-�}ت���9o�L����'�ꍟ�&?bLO`c�OS���Xh��ENFJ��a�ܓتZ*�L��^�������"���${���� ���|�޷ʰ9��#^3���k�Na�CJ��~>[J.�(�k9�m�Xw
��ԥإ^O��NnNe�����1��.�%m�(q*��]V����U�FËÖ��*��^t%8���ҿ���i�T
M���(�o�U���v,�,Ä��%]��:��{�mvO��*����9�B@`*�!R��ơ� ��^��1����=�Q�uS@C8��L�J�+e8�44bѸZ��/���*Ǡk�\�������NmuxM�5���
��h�}���]�65aQ��T�E�V��X໎{�"Qd�����w��e.�׋���Pn����=u���Ę�b���c��?��W���3�6�n�CrI�F�$�vA��.�5�����Dԍ�C���ۉ�1dZ��l	6ۣ��{���kuK=Q��¡�Q�/��i0rH\����uv������b6
�g�^�E���4G)�����y����|�@��:d�0�gC�=���Y}nF ��ᷮ���0j����.���Oy\k���;������Q����"+��@�{�Q�v��a�"6aWo���W!�nyŸ��؉ �x^�=��.z
A{��� �����zJ��V����,ϫq�Q�V�h�hgМ��\xZ�P�&mF����9�q2�H�rQ�!��oY���2.1�l�23���cB����v����+��Q_��`�S ��\����;��{��~�7���z$Md`�*N�	�F2wLژR����c�g�4��K�}�����h<s^�
Nr9E	�VF�0B��	L��Ὲ>�I�{��NMQ�/�D�t��˾�@e9ڏ���v�
�8C�-�2�7e�l����o�xN��Բ^��C���$��H]��\J�5�x�o��@9�,�w�ɗ�I�">���:�� h��q��.�gbO�Z���3>�٪�%��n��Q-������ң��;ɮ�ʋG�!�mԜAb�Y?�^�4"&Z�O%*��?&h˥m�n3��z��'��D��� ���6A_�J$��'����_��;��E����Յ+���?�o����'�Ƭ>�D�e��fv�[�����Ԏ�|1h܍{�����ySw��&�p��=L�vJK�]ۿ��+5nH�T�r����#S�[){�&!NfD���9Y�:b�#��=s#����C� �wl7�E��vĎvd!����w` ��>�������E�9�B9{G�����X�'�⠙�5������N��NEX����=�K�*�����w��1b|��.���1X#BϨ�Y��ڕo�O�г�~��f�(�;��b�:pzLOgª�O"u1�����sl�	��F_-�4q����n�9��(�� w�,-��CȖ�-���O��	�T�b����~��U�!���Յ
:BG�N���q�r��Dv��x�1�>E�;z!~N4�jacE�~5ʦ�T��A�����!s�M�O5���g%MSݷI!Z�j��G� ��O��K����Z!8O@&�'��G��3bQO˱0K��R+(�^�?` 	����u��+Foݱ��1�ոp�xV�$ɜ6^ \�q��3S��n�E�Q-�	�I0�m3�RR��..�k����ǻ��wa&!�pC����T���t.UU]�W�]˸N�S��ݟJ4�ߑ�"p�6�Ч&���fn�K�-Sϸ�^��j'�i���*&���e)n9�x��h�XzА��-�ᄮ�-5�1v"� ��8� ��Q��K-���v�=.>�6y�*r�4�����͈	W��S�Z�.���m�C�L`����Hu�4�������a	~贕F�J��ő�p�k��ܔ�#�t�H}��_+�B7���᫻"��mb�ci����`	�m>�;�쪛�E��F�nQ,\&��q���J�[�1c��x�7��u0�p#���o��g�`Ԥq��}���%�sp��L��9�(��C8�4>��b��
G����Q�FQ1��w�������J��LQM��y9��w̝Z?�z\�����c�3���wsI��0�������wt�3f%ߪa�-{\���2.��*�LQ�����)ke�kc\�wE��T)����v���C�wtY�ύ���vq3�[>���U��r5|@lX�Գ���3�J/�M�[�e70)�����@��D��Sf��(Z�:����ڐ�Q��V%��UiU�z�C��j��R�å[���9I�g����Y�kDК�˚���A�����6r�)Z��b������gIh:;rAү�K�cR⑌L+��ZM���҅���dnE�e��h�`ÇC������G�(�ض���9���}�N�7h��HfD�\G.*rp(�JC쑺��"ZDPS+���9]n�$5Z��s�)���g�	���а� v����H�N��?�b,�[��w���c�/�S�]9ݕ��-��Ywd��a1R��[#96a��"�=r�L���)�,����2��.�M$	E����&(���g�*]!�h�4�>2ƺ�:� �S��Yv�+?>�r�#�� �H�I�Wjg�܄���Y�@�YP���I�s9߱�ik���z�w�
�j�y�a};S�w0���"�i�s�XC>9s�t(?RJ}�Q4�P���n*_�]Q^}my������l�`s*X����w����o���W�ͭ����t�6(��$$7i�*���'���F�A8H�oac�'��5�O2�T��%��lf?!����7�Nm�Ŵ�~@���5&�n]�o�[���-��c�]lE2mJ��MJ3[�59Z��6u�;�����	�l3'4����Y2�h�=9�x�ٶ�=x�D��LTݚ��S������JZ���6z���V���7�F�,��ȍ&���}&�Y��Z��Wy,��2ZX�/TosJY���t*���V9Q�,��y	��%�?��ܺ()�JX('.S#���N(�N�D��OL�2����/��@Y�y����9�U/��yQW�݀�tXi=��f���cX�#�y��3������y=1'���>w��Y�f͍ �n��^K��Ţ� ��n�*�s?"=���h��\;?l�^�"�c��L����S�z8	��y.kO�/&֌o�g ;��9�?c�q"�p-q_�Ȼ;H�,�	�b����,\�29�a��Y�o�SL5�K�#70d���	?�5�	(�Ͼ��4F���X�����Bs���T�qo�Q���I�Z�0ah|�TH;�;=!��S"i�5�7��e3c裯�>�׎\��L�k�~Q���|W6��Q�XZ�R�z�������E�L��S��}ϟqfj��#�'�7�u�@�%���;S�27����'�]����G��Z�|��^9|4-�9��}U�5�)^ڳ���1�>%Oď��pj<����Ȱ>D�q[���XF�Nj��F����'��D��ǒ2X��lS-\ap�Z�4��c�*�d�".&��g�|�Q6���	���&L�r� ��u�J4�\�F�����k�>zHF���}'*�C�Z���s��j ���CJm��7�^c�]�Ec��Buc��f���AA.qwt@�~�r/�8�L�� ��p�=���Z�];�8�9�!��IwսT*������<'ӁauGn���mD���~*�UQ�0��������2vMv��6�F��4.��y��,q���e]_�*�:
����>�l�j��O<9ǔA�s0̨�'��`65E����)�6l�M���
 c" +���R�aM�aj�j*�A��h�վ��u�,�rݚs_�넚�?�.��f*dm�A�!��.5~ޠI=�]F���%^�˖yo��4�3�K ���ۨ�sK�i��� ��x-#ҬB�E����������A@���ں�!��2��f	����-^�߹��l,�~.o���^��z�ecNK@&}7�ĉ�.��򤆝�6���Tȝe&O�(l�W�6�q擥��G�~R�����Hށ��ŲO,L�5�0������s�oUS����|�"�{�â�0>�<aU��9^���v\q�؁����@c����*�Ah�S�Ew��}�s���eV��'q	i���S��0Ե������o���P�GhG�lSܭ� �$wq�������4z&V%�;�6h�=b�BkF���jLY�]N,��#C��H���d:�Bvʛ�)�xs�&�V�}��U����8.��.R��8�%�t�	hD�����I�IJ/cO�b��i`�7L����:���C������Z��)G���F����8Ќ���M�X^�Î-~_j��V#c7�d)�s�����@��U�6x�����B'P�v��Q���L�n�=;�?B $Hd��H1��x����E?�-C�!&���$����*��<%��Y'54�a��/�[�G���A�Y����H��ߡ���ba1\8���K=rɶN��&���*m.���=?��|o�C��X=Z'���_!�;�$^��5���SJxgU�3;�D\�^���iKT������	�3h��f.�#�*|�w<���@��(U�q��| �R(cG�*���|��P<�2K�2����%N��3I!�z�(�GD�&��w@s��~���BA��(��1}�W#�uR�>c�(��̤���%oͰJ�E����v\�[�᫶�x��h�(�n�{y-XR��X�.]�93[DE��^^L"X��)�"�>�_]�┯�s��;�ܖ�(A�=��܀vm?���!\��p80�u�sN�/��
�������#��@j�qz�tŻ�Ə�-@�C�p'A����6��l��^�`5Br�Or6v����g.Z���M�m�xK�g����\24�Pg����00"�P|�T�خ��y�<�'P�%x���gR�FuTAFkh�P��]�A��oL$�NŇ�t-S	s�sRnƠ"�ABĢ�_IԶ�m*��"JX߂I�W��.r��R�6�tG{OWD-C�'��.��+�=�����$����ཋ�ύ�4]�]��P����Q����{W��Û�ě�(NF	}GU�f	C��wO
G�}���o�	-DUs���zH�oʀ#�ț�'{& v��jח�d+�(�p�.6��RIM�D����f�1��%�S0������& ��G�Đ�A�\o��ע)�=����:��a(!=�t|��؉.u ���E���Bm�c�¬#ʵܨ7�ݖ��b�nB�#�L���樂�a��uj9��6�<O��B� Z���Kzp��ų�D��Ý���W� �C��	���j��r6Zg�E�^k�-�&��\k��Kd���aw��6���1D��ht8S"�lީ^'�:�HX$�kB��(�a����Q��p�WᲸ&�M���W!�hÕ��H��������;]>��S�7�G�\��%n���U��k�M����)y�B���� ��p���3 �$�a<��V�!�����;U.�8�����[%�k~d���%�Q;xo�����g�X>���lX�	�����[����!�q]�"�y`��|a)���{$����-qƝh�����8U,4����\��B����\���GP�墂�V���K���i�*�R\�eD��e]�p����԰���� ���tu����[��d#�Z4��!�e߃9��45��>�'n)ɟ���������䉉���ݕ��kwmv\X�O��-[�_��7cRY���d=��	�dg�Ը%�c��`����#65Ld�J�Ϗ��l�g�lŖ����8����4�'Cӕp��k�%���$Ҕ��{�[q�
Ho�G�����5Z�2j2u����o.&�R,m͚H������q�u�/���Q�1���9JI����D_L	g�X����5!��A��ʲu*��l������V������!�G���*���5C��Ab�o�Bv
�3�Bd�j[u��9εT���+�3��&h���P�"J������#c�@J���T�O�AM&�/ͩ'~�b��*�_E����+	j[�e}��'�ɘ���]R��6.6�a�qJ�*�7���6��D~��`�qs�/�M��D1��������Ɩ�ي묿��^E�5̆׀x��Xe�fQ�A�x�(YUXeAU�.�^&cU��M���o��~��Ϝw+�ˀw�\�,S'����=���a�X��Á�&�\���*��hK^af��}�cچ�����A��xM���Ů�n���y����S,�.p��(��1���
٘,�n������i��;�pһ��Ze`\�)�%��Mֈ� ~d��&���P��<D�0�qT��!C��C��\���&H�w�a+ࡶ��"w�z���DX�?��:u�_����S�*DC�D��La��(o��縕������!��������N����+�1�S�S�P����3�9�(����il���gP���sq
]�=��Y_�����~?�z�o	���q'��^V}�xz���~=z��)�H���V�Ws4Q��O�:!
��]�v�������#��5��S���Y@������V���B�_��Ok������	~r���Ja��=�X��mì�ǿ��S�"$aME�BpW�N)�*@f�W��QǾ
Lu񚜝+c6\	�R����V"��9�f�S	�Ar�z���@�Xi(Pu������ZJ`p?4	܏��VDg+���EC�C��\!K�;����� ���E#�)��|����h>��$1E���KК��i!���&n^ b臔��`J�0�������ƅ��s�|����M�ȣt�հ��ZnȬ����&�R� �b�~4;x�UH�;�jǆ E;Y���j"+��^A��%�m�T�]������S�kP����/�H���4������/-��G���O�̉�׈���3V9�%di�o7���ұ!+�Y'�#�I
� VF(4�Y`�G�L	B ?�sDO@l1��㘧j���J�l�����ڼ���͏^�ߕ"=���B�FtTT�[��0�2����2�`��?z���T��|�OLDދ�%�I�����<��W�'�l���	_�.�ʖ��+�j�-���8���ed�؉2D�@�iN����Lr�|sX��](�Cχ�6#-�D�B�1K@ڪB6���=O߷}���;��Ӗ�Վ߱��|�a� �D���q�3��1:�LC���Z������(Նݗ�[��D���A_��0��g[=��y��̀��/Z�l@��Uw�7�ʦ�N�^吓�s3L�u�'�_@=N¨�b�l"f֎pt�!�l�}v,�/��=�%2E#�!t8�1�S�~,��>�#?5�&a>���s	��f^��h�%��,"��9UM�7f8|��RÅ����o��%J6y��<q�L�G�dg۪�ŨR��X����,,�,����\�XWְ8G0���S_6���b�G\�xי��1*��'�U���9F�-��4
㭂��M������f|{��a�sg>�0 @�M5���1_\��J�n�ժOj��K�{��:ǈZ9R�B���]%<[����UP����"�S��#�df!��
�&%� ���?�N�xQ8�g���F�c�6��7m����)���)T�d8�n�J�y ��4�Ҽ<C��'.�Re$Ds��3�τj+=�!-q���j��ҵ �*�Nxz��\$����F���$��_�Z���%�t�k&��ql�����b�F�������AG��ƙoq�6)�%���]6�)B�@`p� o����D�}�C�\�Cծ� P4�]󖆡N���C�J�Y�)���~�uVk�)��{3���Q����$��Os��
u��c�@G��x5����X�]�KS_��CC���kא&p�r����ƒ�}Ւpl����f9�!��)�]����RN��o2]@^+�icm�2�V�r�ɔ�6��d���Yص�h���d����t�m�>���r �ڳ>U2�x���bKt�M4m�!R�j)9hA�+`(h�T-�[�7b|��n���V�7y��g{귫�r_�ʺ���������+R��#-̫�*~8 �]��N��J��v6V\䕃ej�4�GC�׬�T�d�"y�s`�_��.���1�hv���N��R��j:�n�J���z�t#E�N}m��
��B���$�~[���V<�3�|7@���@�WpBO���rׅ��{c���~��D�qnd�/��SDiA�0��J�y�\�������IdB��I��9�@S�!���°���Z���CĀ��&&6��?�q�ˏ��A��sm����}�c9����B!�+��#���]veVS��9��`�CˣТ3[�F�C�a��~�4��Kҡe���������X�/Q�V��e��YYz3s�XK��9;k��'x�슓^�}�"�ѱ08R&������󉧪��K�D�D����
�=�f�N�������McP���Jp�4{���^_�F�2�}����
�!��V	d&��D��9 A7����Te;�_����E��:s��'n�	ߙ�B4a>�k������p�nP�>�n�~qw��Ʋ�T�u��l�[Z��Rm���6<h��NL�a���y?�>��%�f�#����bS/�WL��{Cl���m*v;��� l���Bg����*��\���p
j�5�6OFW��[�0x�o[�()]_�����۱;a�������y�E�;��l��)�q� hb2oʭ�j�������7��顉�b�A$�-k �k4�t���Y@.s���9���	5�w�wE!H���$%IԤ�Os�¯&�v� Y_���u��S�;����+��x���?`�r0�q��pR�uq*`��:��a���9y�E�b��l��62k ��}4�j9��q�3p�����Y=�XRXn	�Hl�nv��?���%�5��E�{����nt7Ue��5L+KG.c�M����3�̲���l2x��֗ض��lD�~:��Z���JݸH�^�m�ǩ�\�B(k�G����I�_V ��� <��OT������C�K^��h�Ŝ�˕*!����|�p*j�jp��Zj�����GǸ�}/����3p�2����1�7��;��0;�[���O�`J��}_��X���ǹ��� {���R�+8 b� �@�ɞBS�b���/��#
���q�D�3��@.�w�A+S�f/}p��7�����x�6/���-LHm�G�u7�b�z #���/�(��<��,0��=�/��]���hc")��W�R2�Xr��x�@�@���y�9��w�*��w�R���E�.�]'Oƣ��V�+u�'��+�cq�?���0�A��<����0�# �nO+/Ǿ�R�1o�e���<W�7��:�?��_q0��.�~��B>��_u=���ޝ����E���{�v����`
�V!��a!E "��Dr,Iz��o-|-��i�:�k^CPS^�8�+����r����q��w��5�FejD�7\d�р��˗̸��1���C�����'���Ov���`{����M�&�WE�.�CG������t����&��b��{+P(s���ᚬ�`����HC!��@̵�L1}�#����u߫�al��&��5Qn�gǿ�Y+�. 5{��`��^}9Ry��;xM^����w|(Q4��YBR���A�yg49�#|4W<�b����h��k+w�A}p�Nf�g!��EL2+��$uC����YW
��2��4�����!I�UAՅ���Z��S	�R�Y�qv)��yj	7��/e�������5�#d�T���Ⅼ4�]2��^&�;�B��� ��`\r������ƧޒX���gƮ�ml?�Y��(���1�Ȏ&ۄ>���� I �A��M�9%�/�
׍W\V�x!Ah$|O��ΜA���XI����!B'$CPP�Sv���O��5_���W	2�`ݟ��B'����c���ԟ#i��<Bo�,�֩h�yp����1gپ���3�e��Q��G��M���au�����sIa:��j�0F.�]�l:�Si�T��`���%��W=�@�uGk�oy���	d`/ (H�+�
p ���&�W��%R&�D
'
Ӛ��8��T���\y����h��=gQ�����5���Ic^�3P	�����&��h>q@�$��7���fj��P�NDhP�����ID�$�4�r	�ղF;J���ט
:�8�8m��*�n�Y�=hvjv�̥r�����sn5�.4�v�"h�2!PD�T��Ɩ%���a������5ˤ���b3uE]������H���\���<e�;�I�a�lgK]�2�*Z��3%_7eHk�:��O��F|�I�f\ft��~�,��z�/���e����*Ās#)�k���Ï`��PYXQ&�۰�$9_�%���{����ܼ���1�BrO��1i[Z))�Wd��ĳ�;PWg�ri4����v��� ͹����8C-���L����rd,��6d�g+�/5�o�9O��P�2�hr';�G�V�?�7Y�k$q_�X�fχ�{_����_oJH�eZlz�iB��:��`�	�t�(�d���}㣶	�a�N��?�Tn������<EK�n/��;��e���w<��3�u����n�a��O3��}�u��: C�� M�.A���\1��%ғ�"-�C�NlH��Y\ֱ"��i�k%��<�q�j�_�헊�n¼r��G`�c��Qj��E�����V�o[����*���H�D���-ae}�h����'��0�9�M[������Fe���Y2�k�0�~���㕲������Ҟ9��BNm��yBp���P�d&7�b�߃���W��ĝ�� >�Z�BU�F�o�;�W0`������1�xZ��h���
g+�@o��?[S�����<��x<�zVflU���5`s�G�ښ�\��N9�YL�&�&}߇�RZ�%���r�g"n:a�	�����$�	Kp=Fh��PF�,b��Ḁ�s�ו����JK�(�BR��'�4�Ht����f��^AX�N8��	q�����1��Q�j�r�j��//��A��N�b�[�^|�MF����Q���2�j�P�>���r[H\��Es�磑�����#HV<�!�l����}�����يuՔ�9�����	̐���"����W���_�!��?�Ǘj<��F|���J�t�>�@���L�7nR��F�J�M�!58�*3%:Tبom���Q� -N�z����ո�`���2)~���UH1ё�ڷ��^�,��w��J3O��s����W���E�0�:<�5��1/0�ύ�`��<��4o1wG��4��lj�2��+��x��`!���)̝�u2}����4��g�/Z{Q�+í7!�o4br�����WTV�A��ٸ9Ɏ����Ñ��;��m�Td~�+�� �W�I��c���6%6xj�最.+�O�`��������\~,�Z��÷�4��		�<�{��׫�z�(�7\�s1��v@	�{7G�y��mf^��/}gJ�BΖ��w����"�+���z5�D_X1�{�r=>��]P[�����]�d��v m����\p��`�.�� ?�Zz��0+�YJk}߹k�����d�T��xn��L�5�XQl^��
^��ȹ�R�1!k��_������S�������g�u���^a���A~�8	_���B�b2ĥ�����0��#�ã�j�-c�F�I���A�͉3���7�l�T{�S��/�<	�d}餅\%MG��J�DS*w�Q��@;E�;dQ�F��e�ww�<�����2�L��gg1�7���>�92lH~nIe�]����¯��T�j�y���(V�ʃP��4|_����Ϯ$����;2	����~\d���g/5��`	���$SYXg�'��$Vϐ��z����K����`Cy&Ow\XD�T��{���+�#��>�c{�U���Ʉ���
�J��W�6��Q�7	6&�Tӳj�?N6̫�K�Ԍ�i�K~�~'#�%��{`7e�#�X�8�qFί�>�' y�n�:?�Y�sO�d9�����#��-�e8v��J�0��RyKT^���a�;�̖$�!�"�|�6�k�Ӡ�Y޼C`�"�ڳ�j0��DƜG?¹7�5�2&wh\8�D���*���q�^��s��?���Ex����y���AwJ�o����VUOf�KȨQ̟jh����G��\�:��w�ۙ(נ��}b����B��}�b�?�'%i#��p���ֵ�y?�z�v� �cG�(��ܫ�J׸�3�&l��}��������/a�v�:_Y�/��MA���
��_��$�����M�T#z��+s�=��=�,�|���l�6��i�O{l���/zMq�8���;Y���
�s��,��Z�e-�G|tN)�/�m��a1m�A�m��Ɲ�����=�_N�� �!g ��w�TF���r\� k%H�6�hc�F�C����g��,CA,&HKx@���L������4MsY����u�P��9.�ncpY)[��83Ѓd.�dĉ/4ʛ2�]D:��e�'��K^1��>>T��+*$�LV���8�j��O%�;/&!�������:P$��t��_M��wN �J�,\�=��M�M���|�48^z��1�5`u]�a�����"]�Ƒb�^G����a�����6�#��Ot�5�]5̺o���[�l�ry��2�qz���F�����t�[#��D�����L咈�n��.�k1^j:"�}�Ș/bΌH�qOa�t-����xw�LP}����N�)8�r4��Ʊ^�c��7��<./"0(����'�<�bm�4o�w�1忧o��Ģ����a�33[
/��I�!��ذ�M�ʩL�~������b�kxbѐG�7m�^5h4�]�b4>n�P�0/9�2���\AJ���𒈐�{��B� ��6꘯d���jt-��B�}������3To�U�mQ�5	 Ek����Q�_�x����3d�پ�k"�_8�iB���cP�dhd�Ú��9���i%@'"�F����ܰ�Usֹ|F�ē��p��^�5I]W��Yh6�`Rg#!�c����fn��j��2��͢W��َ��2�4�,�G�%�+y����B����/U���w�Ťd>Yb�~w���%���|��бl.W����ow� �h��kx?W	h3bÚ��Z��< f�Eo�pz���[ɷK��B� ��9tQJ/�;t��)�=�ԥ���X�RR kϑ �Wm�k<�l������`�]*�Ś��Wd��bB���h������H��c�-�P�������	ɛ����j]	<۪��Mr���2�$�ݴ���>�b�|_�ΐdQ�$���
+����(��Pr?�E�<��{2A�.�0�ߟ������e
�\��F�%�[L��V9�����y	1��2����q�b��:�G�>n� ��;`.(���u��L���c΃�j���#�y&�����﮳�x�`/�LkE�MT�.�����yT& 0�yP�3��]�f������"�7�V�p(j�-B���3ƺk�}�
�/�{��?��V���i� �j�3V��kV�l���x�R{M��& �Y%>�i Q��z����K>>��~���R�KX4(�x�_�媡�qԃy��ݽ��e��IW�;�N>n�Sl�bd$�q�='}M�Z:�Ti�FUv3Ig���'\�2y!�GzN��W2�s�Û"���j ��v�N?+P�r|���\;��R�J'�/�Sɝ
u�Ƒ���f��c��gga�w�=� n�xA�A5n��.�q2�����'d�/~���>(.ǢT�W�$���oS-�L/X2 5�?��.|���#���F��� �fT�޶*���(�W)��(Y�9T��=.�����CnW\���g�)C���]���<���%�P̃�=|�{��e��v7`/_��2�q�X�5{�~l�j�TI@��߶���>���n�����M�B�:b�!K����/�.�/���J;�U3�h��{L=ǃ�\<g���K`����,�o�]���*��[�d��;�S>���e������LC�/�ҾPxo-z��T
[���ŀq����]�8ytqB��9gxC9�e���n�l����2hv��*3O�p�ENi�$O��z# �3�3��$�K��Ő���V�F�=�澼��d~��^�л��q�ΡuGcb�/\����u��l��#���t%zS���iI�z�>ڤ��v(�pP�Cc�t�x��%� �� ��/Q,}�i�ו�#.���
�_�Q�|#�y�~9[�l���V��Ӥ^ߌ����S��@�S�'YkM� �q�ɸ��O�'ɦP�QF&�JQ#�Σ1��b��&s�P�a�[��#�Uhd��B���;��c��HQ6�)�Oywtw��(ϋ�;[[���P\`#^J�x��m����[�Nvs�ܹ*~�MI��ݖ|��5t!����,6.�/�$QB���#��wJ��yPMz�:C��(d�1�(��?~�V��4�dST+�&���M�����ڈ�q�Mڊ񠗉��_��0�bI��I��`P��4>���ui^N��:WՋ�"���(!���1��X��-ǔ{����M�P�%[��.*�S�;v4}�)����-~��K� ~J^r:�}o���1����8�A�ζBYoΌ����[=P�>�Y�C�wꑚ�f1/�ߒ��f�2�ҽ�Go����H��W�_HY�Fk�=LK�4��6��){�L���P1�Z�-6u���{�S�Î�jct7B��֓i��e���h���D\Ώ�"9�GՃ��Ƙj=Gc�\�c�F/j��{b�ZN�����=��$�h�d�TO���#˝�� �2.[ZK�p���w
S7��I�K�!�ݑ���t�9u�OZl���;���)�.­@껏�8ޕJc!~5dfzhnz�a�;u6�k����	�P��j�x��^���qX��� IT\M��`��׉��HA��(����cƺSߐDZx��dT��ke5���v�W�����m����6�w� ���:m�>�;��� lEX�J�6Xk��#��g���<�z��,'��`ƌU �����Uz�e��9�����Iz��"3�/�qūo-i�Zˌ�L�|R�~bB-����M��~���[?}��9&��"=0����KZ�%Nj���ː�/>�j�Gs�tKT2�{�G�i����9��$���`,:o:C���(a�g2^�v��g v�.��b�ᬃ�}An(��Y�kQ���Z�U]	9���p����l9Gw�%f��$7Sܢ�M��E+��4�=���
��Q{��O��ǵ��d$���� ��6M��[����!���b���k�	�����X͆�h�r��.��Cb,�Ĝ_�O���O�1�uk��y�a�c�L����o�+F�Z��'~�x}Yx*4���S��M�(��}߼�\�U�����g��X����o�C�>�+eu�L9�W��l�@�T��s{�D�]Z)�ԳI�0y;���҃=_;�*P���C,C�l�>��!(]����_�E�B/f�Bqsa�T� 繵�R_H�_1����k��j'^��H?�Th����d�#f�I�w$�?l#�-�+��~ ��[�b��^[qI��e.w��%��҃�޾X��Ԯ�h��'��A��~�a� ��6�WUUacor:ĝ<FcDPB�r�T`x�ft$*d�'V����y,�f��{�B.��ק�[���M�F�؜�`D�����x�n�����͆��l�--��<�+�|&�ϑ)�[�j�����A�#�lӱ)작���q!8sP��
����u0�҆�#��v��k��\�H���tÞ
Ni�<��:�Wc�[�h���1�E���bd*!-/�OU�����<s H�*����Fj��'j�Hc�>���]C-�LVˤ�+݁��ӃR�ۿ\�K��q`.%z"?{�����5�脑���É����Ճ>F���Ʋ9�:U��Y�y)HWW�6�#QJ��ۆ3��Ql�C��1�_u���G�6
P�C�C�%i�*�/���Ņu�\�"I:X��� 7.��Ý�J/Q�o�� e'�L-&���:b�v���M�Ъ��X�G-�N4��mۑi�[cH�$��뇚?��E@��%aT�ٷ�R&rU��/��O���dR|4�FPg@nX�7��u�ҋb]����nld��"��S�S�x�=}PE�q�/�(�L�\�k�t�P���,#Kn��=9�(n7��m��G��Ll���3�������PÀ��ck�$���lKC���?t/�Z����C7�V�N�NE�P%�O�����:����E��J%QS�;�b�],B�½�c�@}ox@��V��lH��m-u/�>�$L|��3� ���n��F&;QH�Mq�D��ГL��8�\��o<�b��U���t:��B�5h1�����qY���o�w��ܯ<���}����7��c�$�Jkۂ�DPF=�}v:��&Z��v/�M}zE��<M_9G�!y�Vb!��Ԗ%L����^���d�K�3	�1:j��-4�(�Ƌ*����+s��${�2�	G�c��xB1tq�(��5f��NӜ�L1k]�{�Ϻq%g<y ��yA�7�Zp2���d�+O��>��љny��k�WY�Sw����Q�.O�lQ�nS`�%�078t�!�.j�m�1=}E*�PƤ�W�@�������u�g��Ύ���8I�RA��d��7�-�p$�a1������ߤ�x쉷O��f�a���Ӵ��|�g��v��ݽgq�x�	�i�;X��s�i�o-�I�W�D�p�[0�*8����6eK��auy*8�L)�3w� )��N`����	 ͸ҳ%0(t�+N�C��B�����&�u�Ѳ;�Зvk���Ȇ%L0�8Ì�����2�!����|<�[����ѐ#Y�D�K��\�ݟ�|���(rA�Qz�KJ���/U�s㪍�{�>6�ļ�T�Y�����C�%?\��Z�@)܇5��?���J�7BL�ȋ��A"0�=�`���Hv�`��3����	T�u+q��Y��X�:�+񈜵NQ�B��.R��U��#�@IK�oˏٚ��Km�:_Q�;�Hu���x
=��?�Z|�crGU[_F�W/TT����W����R�ft���ƋnQ�_M|g��/�*R��?CDޑ����wGcy�ƈC����>�V����j;���r�-(PŰʶ��#�`���r�����Z'dx �-j�"*!�YW4-��A+�ۍ������h���8��-�5`c����'a��
],PMi�p<_�llHIz}��G����4��хeD�9Z�:��1B`I�he}ER��)��� �;����-���~�N[N�Q��|p��h��.����n���2F�m��֎�р��\�瓒
7�
��&�2���u�����U�yK��~�51&ӓbJB
�<�M縬�JKʩ�x�����j;}�ʞ]C��n�͆
�5s�0�Lcm�=�[�������b-"{F�@��;�����T�la��?��@�.	Q?��k�2�[(��Ȫ����R��o�&pv�?�:M�e�U�147�' �L�r���6�B]��g'�:�$�H����X�0�Y.����v�(��}n�Q�=a����X?.}g��������bd-
�MT���F:@sT 	�sM��Ҟ4�D���%�=��
/�FJD#�Ů�ג �U��a�wA�z9p���/	AM�&���X�V=�7�d��\g��!�S*k�a(bo�/N��+����Ɩs��\l}ϳ:�r#EhH�i{G�_C��� �5�Y�� �tjGi5+}�����u!t�� ɴ"'V~��K�c���Mq`N�`�34.2���=��W%�ۖ*�و >���Ԅ������%�f��j/�,D��>p��h�����;/υ���p.��<Tք��Fj�����T��x �c��f,��5V[��J��٨Xoe�vǐ��˅�T�M��]奡y5�b����Ժ��e)_x��qN-�r��� Օ�Mb�U9�e@�k�֖Di����<Ik��X�cE�¦,��g�
m���y�l|bkJ,��|�/8ٳ��/��l�SI���G����iM�6��L��[�w.��epk��K��H=N�|g�J��D��g.&�ْ���7�B�����ø%~�hh'Tӭ�����a�my6��1�4�י�l�Ҙ�6K^[���Xҿ�U�$���g�]?��J����R��Y���W�E���?�sL8{���0�pOO������\��3}�	��C�(������N�����Uwʘ�j,y ���������xf�Y�̂��ᱩk9�N�PAǀbk�K��?����@vJZ���+&传R]3��H��Y�H�;
� ��:�<��|���������S?t�������4qZ[NvSR��Q(��}�`��-O&}i�e��*��7�p"M�
�c5��Et"�S�Y~�l剓�����'���\���_p� �qB�A�,3
�9�@�mB!$g��6qh��BQ{��Bti���Ҥ��a�������aB9����<�=MLl�%p��[�W>)F�"��J�H*�h&���h�Kq���J���k����D��$���ѴX���� "�F��������M��\����4Mݬ��lm�9�)/���8��NIe�,���I�S�!M�8qSC9Leo���b��h7	�&�܁dA2�5w�Я��c3��CPnM��+U~5g)�WE����_�.)���NJ5�3�l*�Vt^��xN
`�*����9g��+�g���ӱ��ox���7�@ )����c�Js��
� �c����Ot�[1��<V�|CB�Rs���x@���O�XJO������0��=@Pb3K�˟��(yF���;б�Ur���p��
y��(�h�9C��No���.�O(RQӎ���יv���%
�'̝P���} ��o	8�N繶�����V�E��8F�x@��{M�U��AE�*�
�bW��gR��<��R���O8JȦe��+�Y�|0źF7��~Q)oWb�
��-P���a�[�&�^VnY5	>�Mu�٪!�kBV��?w�����Ӗ�l���������V*y��f�+9v~ߑ*�0�Mn^�Gȗ��%��E��H�JJ'��g��\�PQb�qL���sLހ+cA�<eW��}����B��|��X�CԌP�����1�y�ʴi����.�{��7 ��Yd�?*(�P]����r�֫ȇp�&�1q���@�n� �m��֓���)VG=>EGUn�I�����b�b�%˖���J
@i�C���(�� 컓0��==����j��C��fB�� Mc�Ң����ꈁ�tH��/��gڦ2�G�WѨ/�OȨ<o\�!��ܽͳmS; �C���/��3�Ӱ�cۻ�]*�2}kY֌�:���t�kp�k:�L�x4�
�1�a�4Ec��+,C���2�왣�O���<Su�@L��=A-D�
<���W�Mm\}>��##ܽ�O]���눼���z]�����e*�|�]�)5��KV�c����_R�2'r�.����j�V=�fT��o�Ó��چ�$�9���<�ۇi:�,&��F_9��$��{�X�A��!��:զB]���g�ʝ�-�ǹ��Ie�˳(����ҽY[�*��e��'�idI�Q�h�/�$i)�� �4���x�Ak����{����k�A3M/�C�b�קU�\}r��EF"
е��K�����'W��h4�r|O�^E�����7��B�����#W����������>����q�v�ַ� |<pH3���/9#&aY�g����Dt�g��! 	�����9� ��n�I�`cd�%Jy\�����y�L4��jo�/����<�Fb0��(��@nwѺ�r	�� �l_l�$9��.��i<�o�� x8�y�[Meq��j�4�0f���D���׽�����)�I"(&쩛�P��c����)��ܑ7�E����=�g g^�'B:ٕR��7P&�&���.� R}7w��WJ���G�_<�+����T����:��l�\ct��є<8y��V��y����'��v) \���xGp�䱩
���V�	�62V�S(~�B�\Ƅ=V�	�L�uY~��)��,�m���t��#i
�~��vϳ;B�9�(�1�C��%��>	���HL�:bwpAx�D-bB�Eѯ	�r���rwn�1��,/oR_�E���u�����]�	vq��Ϙp	p_#���=�f��c���|u9n�[>m��ln;�}�����(i;$U�I��]��{r.ϓ���7�ʯy����
�قW:�F{n��\�F�[=��W���|8"�G��;+.߾�DN_׸���
����&�Zn�]Y�;2���C��ue��<D���&������ҁ�oa!�i���n?���F��.�U!�k�s��r����QD+������%���:�xSx�a2�#���t@��Y�f�)��B�c�#��Ȝ5�h5���>\�I�f�����Q���ʥ�q	���`�w�hIz�_��/┻�S9g����Jꇫ*5:���r�Q��B���@�c�c�H����\����_�F^u�"�(��C�t"y@D��U܃�89���A ��[�ζ͙^���A�}�;z$�R���e�Fo��$��k�3~���CJp�j�GJE>����Z�^�Z�<��bC�L��|<�� �0��
�@��h���=�Y�]��g������)Y���?��'��AcM=Ql6�D2�O[o�뉡�`~~*C��aa��@	~��j�y)��;D����i�;� p)��Z|�A$X/8J]s�去@7��oU�R碈�B,M�&�Z�X"pvCF�o.�:d��F���F)�����J�X��^��>X��d�T�=T���;�{��B����gO��D	���w*�-*}XӰ�uI�}	�%�w��[_zq��k��6nL�����ߗX�Q���;q���ͺ���<����.�:�u"d҇���D�_ph-��F"l-�¨��"RV���ޤ#�픫�����#4~��}b�P��K�`ǜ@i?-=��T(�@а+�]�!T���G'�y�V�(9�����=�+���ٕ3����(�U����Xlf�k<
��{��k�0�`G���қ�SfW1�S��/�^�RI����G�v��V����b�]/��Bجpw�z�B��&8�S�N�g_����bM��v�49c��[���	V���iy���zo�T��s��/�|�jK����A!�[��
��X}�ĉR�HDy�5^�w�T�"�5��T����O}�G��⾵��O1�q��7r����'>�e�[� ܜ|MJ�W/{�W"gAܶl���[\-�s�����R���ϐKpB� �Ϙq.������T ����T`!�y@�*����]��#��q��S�~��S��TW	�~8��)x^�C8�k�'��כIg���6��oz(�}�XΡ�e�S�A��ޓ�g��ɛ��j��7ǝ=�,�|���s.q��Y�>�W����+������>}U���}j��sv�Op��[��Ldv�a��Z
�C��p��|}3Z|��9��-M��M,���{wkx[����	��b���g��"��&~+틉���zj���.�����qf�)R�g/�� y��\�2�����H'/ι����:����n?3)Vp'
����u,0�i���E"C����;J�<U:u���a˜������x^;��
[d��5̶0t#F����l͒�]f�-W�\7'_.:�[���� Y_�V��ݝ�*rÃZrL�z?��ذ��+L��?�X���[J�/��~u\�1<i�g�]��x�Fa�6fTs���3W
y�E�RWj�we� A��@��*"���aG�i#�`!͐Qk$7��,����L$�>V���*6X߈��#���+�����c'!���$�����5��q5Nq����և���t�v0w�Ft[�e�3�fE9�^�����O��������/1���uP,���æ���$���6`;�^� ;OM��W��g�cW�"�uZlDb��H��"\�-����Tg�Vv;q�E˪�(�c�,IA�wE��sY/.P��.26�e���g;_Ì��Z���%�Q�c������`�&��\`��T�FIY9��37��J��2���jv;�7�J!�S�������I��)��43ȜA�������tb�&6�H���  ,���tc����'8%FI�[�Ts������ٴ�{(�q�rxA��fUQ�,�)f�"}�)G���_���?�E�\s^�d*��Ҝ+~!�ר�1��u���cF�4��[��,�8��p���A�د �s�ls՞8x2�A1z�&�ːecd�J���<�����>:��ĆF�K�s��8dΚ[C���rꈩ-;	�]D���;[�1��)�U�����;h(G���S�#�s���3h��Z�V��w�#=0�3r��DeL�������)>�Uо՗��m��կ\*X��e#�1��&�����c�]������k�%	���!u�SP~�-���4�5�j*�$E&	+��q�a�ݯ2��K@��@��@�۝/4ݐ�H��B�H_N'��x���Wmٿ��N�Q�^̝������B���'�\�(H�A�8�2đ��FmWq�D���˹�{�!���G|�A��K�� ��N�'�ѫa^	��)�"��%'8�D���5:vU�NU�Mu6g����iJ�l�#��x:�/ܫ�Th+�-��(kf�_����g8]B䨭#P{e�;�J@���Qv�x���W[,���v�[�:�3�H���?w�Ki�ݠ"�v�AQ�5c��V�MfQ�������~��Yw�M�?�T��Xi�>�5=��0io��=*w��I���W���q�y���^>�_?����BKl�31��;h ���Y0�"K���[����� ��O�_�RR��c\a�!t��k3H}�#�vi�Tٳ>��B�Z3=��3*�Oz�,i���3*�<��@#��ە�!U/�7����� �+\O� �t1NI��ĝ���z~fA��$X��#����|M��
M� �<09
���DH���8�I$�KńEE��F.���T���Rہ�x�.e�̮��96l�� �]�b��%�8È��XM�t3��+���+J�}Ȏ�'�x�1em]��4K$_����\�a׋�mD��K�e:gu7S�f$��Q�3yrEa�8R9G��C��*@�(�<��D�/9A�2
Fd9�b P4h���u�餳�n;[x2&]k���Ǌ����k��o:S����u�@6��R�[DJ��0�9#��7��*$����u6���C��|����M��	Y�x�sX���z����AC�=��?[A�ۄ�`�O�%�J^nJu�2�Gy�l�!��.X���kE�ݮs�����%$5�YΞYf7Ә�tӍ��9�F��/�j���ⵓO�+�_ȧ�B��0枳�o�mF�q��sa�>�d�%� ���ٽ�w��+��|���+�Cb̠�����h�Rx��S}O�qp ���*5��J��=z�$��rG����1:�%�^ط3�6��8���F ��?{���^wC�s�����K����P�0��@ҋ��<6����:�[.�+v��T��K=U��/��,f�˯����h���;���RQdS�ǰ��6/�?y}��X�a⳪+���<*�3���1��Q���Y��%�5�����C��_@��f]�c�j�8�o.W����?��#�Έ,�	����x�E-�Z�x��v�P�3d���1#=��+�p���U��
�F�Z~�L��j?V9���@A)"T��A��/T��!�&R�8r�j��u��kI;�¸².G<��P8k%�a���t��\�؆ ��8��p�bpk�H%�2Q#dhR��Armm���ᐿ�@@/�v��<T���z\�!D�>�T�>�yp�{<�K��&249���ь��F�a�v媒�3�1�ui��/���k�*�b�㨮>�u�E9�q��ac�8;���׹��4���U��>MB; �&�R�\/m��t�G��H�{x�ͪg�=��W�/��̢�ޙ�X���$�6?�fy� �5���.Da�DM��9�|f����[
hY�I�[F�T�T'~1Ȩ\��t�2���
��)5�� �7[r�ǥr�����`!>,�ʒj}e�;���p_ DG�
���]��L�g��C��k�MV~��'QO<������QnU�w���%����H���P"<�H�<�ﳿ�f�����i�0+#lzIa������&�b� �x�1XU��2�Z*��ɶ}���GD�8��䇓��4���3�R��$*cV�(��3��,�B�uɩ���;�CZP�Ya��B�z�4�r��_҅S�}�K�����+6���S�FTz�+7 c�w&H�T���7�>��-B��/g/��x{TB:�q^�m���w�}T�Y�%�La[�&���y��9��F��oz=w�`r�~�7�?|�F�g�2�{�4zꅆ��d��㼔�r���xO.�B�y-qXX��!���������[��%^I,S�Ěa�3�(���~�[c5|WO�(t{�Y��Q:�W1����@��$����;m��υ��i�N���S��+�����|�ˇj�i��T������r�/�����Ԓ�hz�Oj���p���8��R���V#�kC#�%�������a�릒TZ�X�fE���U~�5�:��d����w�S����M��&���:�z@�3�����/%!�R�iG����������ULb}�t�����Yd��23.\����~��U��P�?e��,�h���A��h՘)���|�uM��=�5
v��z���)�9l+~�	n܏��w��QE���J�D��n��tqd��p֬�4in�`� ����Cj�1���mL���=X�"$k�u}�8�����Q`R0�Mƭ�&����q$ȋ	��'V�{nJ�w�AץʙX ����T���˶��K�v����[Az�*�]��#�3����Bq��y˹{�a�A����e�/��Ք��E˦^��Y����[�o�
!��b'?p�0|w��Y^���~'��ʴ�F��<몞�)�Ù�,;�q��0��0��r�
Ә�$m*5�^�ҟl7-_���,W&���[���x�D��O�;.�r��Mm8�sk�w��E3(�ig�װx� t�1d���
NU���J��z�'�|�#�{���S<�Ũ�� �?������5��_�X����̸�yX.O�6���5n�����w�+����|���G�M��C���j"�o�zNu�U�oK���$?�� �\|v�MIa�&�
3o��D�p��{@��P����	7A�w��S&�G\؟O������F��;g���J�ޡ��C`<�r3����=K���e��_��Q�x�����#���Z��+2���!��L��ʜz��8���d�����rM��Rs��ιQ��+
�Dh��K[_>l��n�0��0���(�t�i����&lBL�@"ޗ"��`�3�'�mh ���Ɗ�+R"��1+t��E3����RyE��K�v!.
ךV��0q�9*����+�Y+��C.��=��WC���K]�0�9պSz����=A���p�oê���Z�z �f$7}���Ѱ\i�ZT���5YQ���7CFVC��w7�K�u���q�0�/I	`��y�،�E`�J$k���6�'�}_ �R�1f��:�
��/�f=m|%��/��fg��y/�/_��Sd�Xht�H�Jk{6"�[O*G���8�����=���"�[�#aN��^5�ų(~dz$�B�Q_��N��D��(ӵ6�e	N��8���y��߯
�<�Oy}4����KTQ�@h2��3A�q�$|����_�^gHE~�}����@]����?��B� Fu.r��K�t��%Z��;����GEdV���'��NG��X�C�ь`g{��x/��;�j���T��WU�C�_h7���G����M���v:� 5(�ӥ�,�]�7���,}�&�튬���|��HOWV��%T,�W���@f�`�C�U�����2�GI,ۍt��<LT�v���+!v��Փ�x�mj�G��C�_g#�#`J�]����]������� 0�{2Y!ٚB�c�`�]��}gH9����d����R�OAm+�0'�
�9Q�(8����O4�`�v�����\^ݡ��I&n�����3��&��\��Y@��[.4��=�~� O�YY�73�TOTQ�3g�U.�ڍ?��*K/�~y��~�4��?�/~�I�ʅ�8����g��W/@�4=Bd�Rnv�O��"P,���D�x�N��j��^;�uS�v�
K&�0*�}e��V���CG��CG̮�k&��R֎I��b�|Qߨ~��D0��Nfa�GW\�%�Ǣ;ݙ�����t�c�p¯�$�n���O�>�˸�M����g-V!u��R��x�5�gv����F=װ+5�`�C�w��N��]�q�(&^�@�s�j?���
�̯2�[�
�~?�)Ц�Z�;+��?��0��rS(ʣZ�t��d
�c���Ł�N�@�ƇMg蟛�Lżh��ц��hZ5G�:cB�
70M(�c��Q��wɌl䲺��e���_�y��?x�E#r����4�u��:"��������J9f��s�����|�J�
��bB�ΎÊ�\�����5�(�ꏰ�s�<���ʧ�\���.i�qh���z�v�Z�n|7݂E���e��r|
8����
�9�$�|��GA�/�0L��F�߃�V(K\��B�~���<�ˇ�X�n�B !�&�\ho�ԇ0�)�!lj�t��]i�`�
&�vY�� �_��V�'�{)V�~ܷ԰U��Т�YM�VK�e�f��^!Z]ĖPD����kQmnȥ�em�|R�G87�?���j;O ��ڄwD���Xq�<L�3� �ü�V���df>[��� ��CN[�D�>Q��
�6������_Z�m�D�;&�,���������R'#D��n`�sɪ<ʏ����v_|M��U�.BC�}	�D�����f_]G�TT�ե>W�V 4UF�GgG%�����ǈ�peT�Dr���_��ՎlԤw�F�RZ���/
Z�ϓ�)zH���ރ���FρI�M� cIهoB�.q!���#~�h^��/g��^�8���Ivm'�h˃-~0����p��_�B�
{�G��Zk ��Sh>�(�x�F��:0���z�_#��	�&�Ѵdo�l_��Ԅ3r������<��ʋj]~d���i�5A���϶��ʊjnM�Z�P��i��������h��R_��#����~{�l���J�bE����k����C��xۈ�K[�4��g�D�u]Q�;}f�tgN�U�$RW'��	�+�U�]n[z���o@|�2��:�f�+�V_�nQ��ո�����h��I�v"�LH26��k��Y_%��&p�L�Q����9*!ܤ�RO��T�j��ζ�ڸ������&�Х-s�=5$�	��T6dx�#p��C��-Om�{.4�WL�{p�6�~G��<�&��S�4y��B�ο˿WE�}�P�i�KD^7��#)!�tx�4s�Z;�!R�G*�w�`X�r���ߞIRm:G���;r�#��ֈ'q(~<PS��u@5��Xa�!���z��Ί�U�q^��0��|�1��b�����`����A��?+�b翟���r qLi�� [HC�b�����"��o��ٌQ2cLRۀK�P��v"]�w�T/sg��n�+���KT����� �����y`�E�͌�R�h1y�5lJ~>��Ai�Y(�����V�0l�r�{�
,��D��f͹9Л;�������4�#�TgÌ���&��p �n�U+�h]q-}3[|�$��x0�J��	�:��=�V�Sv�:^�:�5�s@�;��Ax0�W��	�_z$�śp�[���D!K�����}�[c=t7�����z9Fg����H�s�{�8ш޳��UΟ�m����e؏p�ıF���!��@��4"�/߆)A!�������{aH4~N����J6g_��P;N�Kw�2梕s�6~F��R����V����Y�H�@4�Ck03G���]f*QS+*%��(���UOCW*��'{NQb6��[��v��#>4�>��3(:]�����a��A���'��
��=+�����َ��U�J3.��2��04b�Zs��x���N�ZD��{��<+�e)߱���m9���m�?���`JM��DL�㶱
�$��o��c��J�}�1�*b
��<c�8��f:���A3;@���s&�ű�ѣ��_�����Auf���(�˩�����ދFxC�h'ʑ78U���Z5���O��+R"�~'�z	l�Xm�!{�Z��l2v�4 
��٨���:z�te� ��OvZ�7�b]���[+�&
��5q�;��U�<������/���4�o&i�*S�E��o���ᙹV.
��_�>AZ c��?��$kF�ED�����2���J����F��z�n�{6��=�Ae���'څ�i�r]���?�3`c_ۃv�v�8Ͻ��l;U���w/�cGn�Ǯ��Ս	n{L"3I~[sK��^p/��M��	{�p����ہ=������R�(��G��}gi��o���l�Ld�%܄�M�UF�\�_�E�<9��4����}�ܛ	؊1��vhA�˭�[L�����ڇ�r��$��0Q�3c�ӹ��w�/.�F�{�_ٺ[�Ed�񇻓��bب?*�c�{�� ␛)M"��$>�P� h{?�>�㈾��䖉�
��_Ǫ�Uj+�j���$+����E�M��ISχ�c�����U8"vy:�ߔ���I�])�ëŹ�9x�R@�qV�y�42����!�����%�6��)���X"�{ps�s��u�y`�=�VemXjv�k����-���T���qH�P��l����tB�������8�(���y� ��h��>�����X��1,�9\��ɿ�A��N��m�c�ϴD�/������?�^����]�,�o{҃�%�?<\���s$=����Z�uDT��"�)#c��ע�,�i�(Bޮ�8�H=�ݸ{/�0F�ƙ+�[�8V�9��}5�h��c7��E(Uz訂?�yŢdY%���ln$�G0`�B��}��d��4S"׭��@Mr�kv �K ��2�0����;\WH�$/���P��`��3L��<���()?F��xY�
���s�{G��k��0��P9	,҉�T������Z1G`���2m���8�CL7'���ὐBI�����)�!	�k1�;
{�`���F!V��BQ�۔�^�3�9��:����^�V�:�&�� q�S@c��*��͌�|�A>��6sp��ߎ��_�R�m����BLq��3�[U3(@�Z7��.�(�NJ��.3��v�������C��~���7�G?G��董�%1}*���D�@�\����e�*,�7��G�SA�SZ�H�m��&�O��j�9a��yT�x�+�_v���j\ך��U��c���X�_<�R[��p5h��g^H�<Z�i,ru,�}^���]���)<��Cc�0q$��˓�Է3��5i�2<�ɰ2$lA���ݘR�;T��t
Uf���DHC��pq����BK�ڣ�&�P��i��.���ʰ�~'�Bh�#>�^}��y�:��dD-b7��4�l��1�E��Rţ}���Koh��,�vƤ<�NDg���0��e+�?��j��$ō+/�\"�Bas{���ܒ���"��JE�(3ߘ@kߘ�?J�3���a�A��<"���|\�4��	���PҒC�S��d;g���IP��RtGA~��-zͷ��QAUl�k"�e��������wa��u�B������$�������7W��ap��\-3�g�ѭ6����|��R�c%}cӽ��lV ��G�X��#�kN��."��\�A
,=�NA��꭯���W��1�h�܎i�L"�_�2r'�PO'�ϫӼ5��)��}�]i:�
��R�-E�31��)H}�k�bHR�5��	��'�|���S�:�gV�{R7]K-t__x+�q�Ќ6��L������G�ƄmJA���%����Z�%=\��ӒצsM��Z�LgJq�i\�SDd�J�ڕ�|�bP�	��M!鰣�װ���Y�p3��p���W�EQ�:=�:�/���q�yg:�
^�3p�NS�6��Dw�O�N[� S�E�a�s���8�R��z��}ݼ��'���E�"u�=���XR�W�Nӄf��R}�1����41��L� ���1]*�6Sm�Q�պ+��?&���{��]���h��X��,�(�.=Qv4@�� km!d��>��s+�o��X5�|���.%���-��l��ڃ%b�f+�	0Q���dW���)j3UQ�|�j��A��盫od�3�YG�g٧�CLŋ<��|���ףMZ�W��J#��1	JI�n�=�.e��C�Q��G��}/�_� �8S��sx��1f��}�
w�Ny�Z�]�ۘ�x�uS�?�ɣ9���ܧ��$t(��v���hmѷ�6v©�ZP��U5pf��d>�#��[��,�U�J�C6�i�Ű���]��e\
������)�!|H=5��Ɖ�翖C�d�7|ko���/�\nخ2�۠ñl��./b�������j��cB��X����,C/T�_٠e�G�$"q�v��ۙ���E�7�JoUа�5Ps<'N���Fpx�N���(�:a���G�!%$��s'{�R^�Y��}�Hs=� [x�	{�a���s)Ua���N��~�w����}a���aW���8�C�R�����+�B��O���I��k�Twe�iI�٪vI��5�s��I�x�5��vǛ����l�'5�9�]v�9�vB���I���'�����au���9��(�8�]��42ap���d��^��o��jD[@+���^�p?L��_tJIp�4�7gXG�EOⵒ�w�.Dq^3�ӄ}Z�VN��Я�#�tC�)�\�����b�%F�c	Ծյ�p����S��G�!��'W��;��#����f`@s*���C��u���Z�)8���+�%fLQ�ϙV�� 04k�S[�]���؎%����U�s�v�v�!�A�?Sg�Z!6\���xm$6�͉:��')2	�~S�Q+�puF؊r��E��@���{�����a��q�W��$8��.�F1�x�7q��\�f�-�>�R�ͺ��B����]s�)4���Ɔ��[[Ѻ����9��Xw%/}�C�Y��Z��H��z~P6iX�
�|K��~k� ���	V�7�+n8�W5����JP���Z�Gdￅ#�
���`)��V����s�v�#��>�d�/��d�ŨI��og m��*�g1�<"��,��"AG�O,aG��d]�n�	�-����B8I�#�c��MEJ�6���{���'��I��v���v��4X9@T�( �}��b���b��F�3�x7=�(c�ωM�X�f:7���c�����̝�d���A�\-!�W����^£������f߇�x��?u[��
�)�����_d�,+�ձ5�m_hN�HDa���I����U���*�4��Y�7����{T!n�rU	�z'w�;.�<#�W&��ho��s���|\������Y�����*��*���f́EZC�trD��ߒ\m�z
�x���d�R�yo�0s��
����K��HL5�K6u��1���������6۫צ3�a�l���S� 6�c��O����3��MHF�#v+����2�H;���}h��(���9LY�+���B�6�o ���l�c��1#s��Oo���q�/�oA�5ZVd�*l�X"n��7��Y-�L�/Sm�}e��6��<GZ�0�NW7�_��_�_Fa\��KV�gԄ:��ҷ0�_s.��s����5I��]7�N�>y$��H����OT�Ld�,�������]��AG�9p��p�������-���D���0͵�����ד�e�`Ex�2^���1ew���r}O�.�EbC�`a�a>.#�O������D0���܏�>��F
�������T
n�������x��Y7�h�١�B�7slp,��Î�@T���L,�04"me��Q��Ɔ�EW�kW�ړ}5�:��R;@��$� �X��r��+��-^Y]<�#�<��:�b$����.���	O�u��,7���|Ί��ro/��V\Ys��!��\�EZ� �T�}�=E�vW�)����n���G������~x|�gk'O�!�Yt
i�L��K>��G��s_���*�����癟,�M�$-Dd��0�ř�m;�y�pd,��C֐��,�N�
s�+d��0�/�[2M�u���2�"Z=��?ª���XP)��Z��'���mFO^p�&[P����l��t��2Z��a�F-���O�T��-Ҙ�zk0�K��0��v}�U8P,�0��PcTu��׋�D��"�f���O��z}���w���.�w$���`�V k�O�E�1ީz�,�;�A
�x���h���KB�zO����%0��=��3���I��3R� ��F����xNu���w-��2�ȼ1�`��I_�o �ؑkϛ�y�ѕ%�r�mfF@��^���K���E�y4�ry���w��[�����#̂P�������-aV�R�ìf�I0���SٰL��:�8L�-�T�� ��=�iʆ�Yfz1�{�E\h�u�ޟPf)�Qڇ�Q"u��" -l>ߚ%Wdе�����������`W/"��ܠ<ss�WHJHp���{���~�1i�,�)���a��0?��X���h�D.˿)�ʝ1�4��ϟSĥ�f,�>fn-��؃7c��y	wR��{v��x������i:��\ h�I!M5�z��Hyz�z�_^X/�8�T���RL0���՟�2U�����8�pɄ��x� �8��?@�Y���M�l��g ����i��j|E����j$]�4��x�6�R�t�S$'<a>���ś:�~}T�={�Q^��v��]���j����n
��B�b���	���	��G������*/�@=��տi]x���������iAa(����%Qː]�G�Π��,A6q3�ݐ�q[���3��x��&��,��<F����N &￬����%O���,�(�B�g_��8����kq��N2P��V�B�\�}�a�D븨;�ߦA*�����Åv���=¼0OM�"i�󹵃�m�G[.~�2D:����42��9̄iA�'5�J��VW9d{|�`2�^��(/�?n�'�'�v�W�b��I�m�֎���G�ى�v�7��EX�J)�I��+r���B�$28�kt�O�?���i��O ��Ъ+�)Zv��b�4�͌ϲ}hc'��>&K��H���b!���D�{v�n}�$���n`�d�D�Н�O}��	r+<�h�I���2�fK��%�>��t?<��؎=�4a�~�����\�}���/�����d��������i3ѥ��ō t��꬗7�@Vm=�׏o���I���
dG�4�`9�����gUVS�!�����yNW�>%��,�=?�]@4�jZ3�]Ø�/��Y��fmH�٢=�;X�6��1x��Z=��[��_���I�9��p�oyy܂ab��TV���y��Z�r]!�1Ҭ�Ba<�T�2�~TF-\%��y�Xۨ�������O	V�>?Ȱ|!�f?4��e5u����^JB����$��(P=Y�C�Ӛ�S.�f�A�T�>Ⱥ{��]ZF�V;����v;�,�a\hsk��Ɗ�|�umo_u/���%υD��C7�'x��#�>T����G`������o��X���s�	�t/��������;E�u�'��\�3��F��C(s��Dw�HT������ ƺf]��}>��ӡ��qV2��.}a[?�u�`5�Q�
�aq�|��T.� dUSX��k�ȵ��Ss\<�z�SQ[�َ�0̘{k;��:w0���Je��s�h������+�파��I%/cN��e>y�HSsRX�b�Z�{
��\��!]�'i)]Ti�/0�t9X]k�$u��Ptv}i�($%*���yo�y_�&/L(|/��NU�Q�dgun�y���8���Z�-ޜg�|�G'�q�����4� `���X�,�x�]D��K���>�����1�|�&S�Od����c:�̇l*"�ܣ ���
�euH�'� H����2uy��G�ͤ'bJQ��-<�x�̓�>�=��aVWTd��JGR�[밎�-[�N�)���Úl����)��[�\��C�1Z�!;�L���R4���c��h����;x�F�ǡ][ ܄�=�b�Qu���΀��W��F�'a痄��.�(�R`�q^��_�AH��"��g��Uk�~'��Ó�ZO�(��@S��R8�m��~Cj�%�H�p">�F��X/puv'�ܼ��[�A�*����
���!X&T ��C���}�v����t����;ݺ�	�&}���\!�p�pEq��S�������>�������*ݼRB\ �]8�n�]�p[H�Z6��b�;@^�^��t�-�����~�2i/�SQ�����x�X��:��A�����mg���E��y���U�K��\�F���p1�q�/��ô�M�ԉ~Sv6�5<�tIN�4"�f������x���si����O�=�t/�(Z�j�JkOqrD_�FO��x�$�;�3L�-�T�2j?ö�-�A{��$�1ɼ(_.�0�C�\�9m��9揓�L�+�k4���.�����D��_�˓>��j3М����E�����P"%��h�3�b�D�V���[��E�XE��{�_!���|휯�9賟�`NIEI+T�$��d�t�}��VUaڷ7��R�?�l:BWk|��0"URAa���%W��6x��N)o��L�z����i����r؅�D�.���Jp���V�U�F���¤�T#a��b�UX�ͻB��t��kWB����Z'�\i���u��NZ�<|��2*��T,��D��b�����F`���n+�$�s{aE�b�O��$�I��{�T]��YJ��e0~_���-��y2~�آ���$�J��<T\�AV��D�s�W�/�
����w��z���ZI�մbG4ٖ���?���(Ҷѹ�;�۸�w�)�+dǳ�bA���z5Jc�'����YxZZD	Vw�6k�N#�T��L�[׊�J�H@��<h>7�K�I���lz�9���-&�F��rA���2�� ��0+��$�
)�_�'�hu>j�넺��z�sz��EN�PPkI���ЄS�ef��k|�e�.�AA��D�U���R����]a�]))\F;���KK[�xY�pk���&�c��3PCt	>���)%B�����ݬ:Q���� �����r+�\�ƙ����y���~ש(�v��)���c8��۩gw��,tH����%�%R�@,U��Xz�(
�|��#���=o+������b��{��7�3<ë�<���K�{�J���9D��������1���jTx��8h?p��D�ڵ�V7Ș��1�-XoX�b7��`L�^s�-��L�gɜ�;xJ�n������^~� ��a%2����[�G?m�T�u� �v_����߱��B$H�?�B�z���(^���e�5�|d�ó��t�w��S��a�x��~�<�\��m�L+p���<̕�݉�½	~��,��0���r=�9�6�oG�τ���9?�Z-|����\L�@4�=�АR��a�L�=X&$����r�=�z.;~�.�/� m �9ӁC�A�q���΅�Z;ki4J�]�����O���A�H��.8�)9H�N��˙M��5;���D̻R�O���S��o���o��=Hșf�<Nn&c�0�q[��2�� ݸ���'͓U��Li~B�;�o�PZ1�M!?�ar	��C������}N��n��2�@n\�򡜔�t�J?&`f��������vJ�m�Ⱥe��~r>o>KY�p��e3sC�u_�/q�p��'�30����H�	h��+��0�:����]���P>/p��!�����_�-Y����f��hρOH���%^<΃����\q�8��_�7~@GWc�5�<��~Ջ-إ^�E��41�7��&2z��&,���g��n�t�ˏ�ܯBp���^���ъ|�Nʡ�s����c�W�0]�%�<����q�k����X������mB��0�jNds�5����SP����%B�b�hw>`A����Sf!����t��-�{+����}P�b�:�á@��կ���l	�<嵭A�TKB�"��OL���u�t4N��
~�.D�k�#t��hğ�9�����?�T���/}i��������HI����ƍ�%^�
;���~��"��p�Q+��Z�.{��q��~��ρF�Q�{�D,^��l9�=�?�p� ���b�>i����3;���4z
�Qَ �>�0$��<z��Ր׎���/�9��������p�����:o}�>G����#0<^������Dm��T�E��{��*��q ����ld��2���MOW3,HrTү�͌�(&!�-q,�(��Qj����o�����!��Ϟ����_�����>p����?T�=Sك�co}� �M�H}�1��I�Mqpƴ��l�^�]0���>Y��P�q;N�@���0����9�)��C0��@��DQp���Q\��Dϐ�]�+E�-.�[�ѷ�u	�J�7!-���x���A�9

9�u%Sx�,G���xm�� �
;��C:��gXr���aG�6�S����y?��$�sH%�}�]j��T���HՀԘW��D�5��gI��ǝ����l�G���a-l��6-�{j�m>���X�Y�� B����m��I��T9�C����<�H���9+���.����[?�C�w�ˬ&D�8�X��깩�g�W��w!�L��<�)�7���Ϫ����+3�<�#�'8��|�":6ag�>��!-Z�39�j	�w�``k��VyV|b� ����7���(:�Ք	�1ϴ��jɩ��kf3�������g D��/"�H&`%�nO�D����c��'3��;�Wi�ܘY� j�YԀ�q�MU�6�&��/��n��3~�K͐��]�7��y6?b�@v)�3��|è�VF�~kv�D�#�F0���v
7�zE�('P�Jd;��~��-\$C���3,�$�|,kL���w�Az7)<L���i8	h�r�'�±���4���`_�0���qy3�@Md����>l&�N@w��@�Z�-F���� ���Y��yL-ߙi��D ����5��A�dC�k�#�foN@
�P��ii8�Cml4�0��7E�z������^lܿx�ӵ��N��5�pl�`���bx5A]؝�C}��s�u;�b�Q�s¥����Hdz��2& ��j��S@y5
���������D�͊�$�����N��̒�A��!�`y��R�)xx����'�f����� :�"(Pڢ�п��B�!��~�L�\z���Ni�~�=a�Oo���K����;�M�м�q�1G9𮪎r�U���M���m�I�6���딋O@M!JMM��oȖ|=r8<�y����jXǿ��F��7�b�.��ҝP�)�/�T�]O4�B�C���`�(�'�`,��5,���O��,JvdI��B7�fD1�Nڦ4#ΝW��2�b8�xu��f�P�����g��&���T�e��*�V~|�7�&�tA���qA�j����LL�H�w�|M�]{ni�u2�I���zMջQX"�]+�	���IH�_P�H!̂��b����a����>tJ�;�����[L̐��/���&��{z�=�
��O}�F��1����FC�����/�@g T�Du�@܆.�57�_"wa��Y�P~�P����Ij�����PM�?�ML�9�W��&�\��Nǹ2��?tXiә��9>ʽ����܆M_�\H�z5���yЗ�����^֩��4��Up
�߲�K��|M����Q�ϊ�	пce,�k��ٵ��h�V�w�+�R�5�9[�����i�~r�P�1˽��A#MZ<�Ž�O���9Uk��;��!���"��v�F_7G>��Հ�ٿiZ�J��n�Wx-H���AS���v\V�7�:yg:rG�FyX�K韷�n��2�?�ɍ�2N^���E�D���t�(�E�dpx���܅BLX�[� ZԽ�)�L�Y�%�\R���m8(wxK�@�B�ܒ�j�WF�m��'z��`>4ȧ��e����e��^����`�~��ҭ ������G?��(�cP��ʶ�I�D�"�u^����.��#� ����2]I�N�#�C���߾����ڬ+i�*6}M���K�Alg�Iމ1=����N�N�\�^�҈��1/~�n���+13_�w����Oiμ?�ۥz[�@�b��%����2 c8w�f$�_�h{LfM�ޣHHm^I�=_�0�_3�oMd7�Â������&ʶ����Z�=���ҩP������I�j��@%�Z�͹�K�f�,�.9����ޒ���p@�X������X�iɐ��juZ�j�#}����1E,�z�z��2M޺�ZX��l�*=|u��3�@ߢ��	c�ej�_k��Ԓ�.�2
�3�p��'�DK��[�@ml�<���,�w�ht!��O���ٱ%B����Up���ÿ����lt�Ȯ�ԧfö��1ʽ0��(܈Q`wQm�3���U�Bz!��Q� '��=���N��\�"�2� J��6&1xR�e}�WR�k��ӌZg>1����|�ijQVT��/c�yK�.�I[*�\:��`��?R��8�R6��l�����]�)L�l��?R�'r������e;#Y.a�@d՚�eYthO�<�g�u�`��⊧*S��4"�풐�5P�C�<	��(�QBV������b_�Ң2��e�S9'1�i�0��֗v15BY�JJ [E#p^.z Y6O�2�X����^Ӓ�K�Bl�wy��|s0�%�R���%�=N�t��>x��Z��R_q�l��i���\�\ި!̸P�� q��*���S䲵�~m\�1)�Y%D�L����!���k��{��$�>��0[!�	?!0�s��%�^v��� Pc����YNXѳ�ߡ�3��F�|ջa���k=�vp�:M��3_nNG1�E�ś��!\��֮M��M���E�������#S�'�<�oo\(�=�|�e��y�H�n�@�pGy}��f{A�$pİ��@�m� �������r>�"ni���K��8HR��6����@�����}�,��;���1����@T(�����m�0#�9��W�K�tO��@ϲP��AK��.2��+Ӛa�����pio�T?C��-�Io��Q�l��*hn{��7�{�W��9���W{��9Bd�⎑�g�	�O��
�yn��E���gb$`ޕO��F��|�OU������?�?R�����'�.�p�m����g&ȇ1����1�+�X���>FN!��s�}7�)hC�;)���v��0���.�qG��(�M4��>-�R}�.T��9�H��o�c�P�9Dԫ����.v�`�#Z����p[������n`����a*.���W��� ��֊�_(K:E��B6�D�C�N��{��.G�n���Jۡ� y*���^o����U���3��p���n�5kM2袜�6�b�����2�2�b��ڐ.[DDF��I��Y8sZ�\�6iH5�1�������PȨ��Е�5�߷�Ѽ��EW�[p$q9����[!�~� �Z�t缺A2<`iH�]s4v��W:ڃTt/�=QEJ>���%׏�vJ�N}g�55d!�gj�̾��b��	<./���Wh:>����!�-2(�� �f|\�W.�K��@t�2}�\^����.�e�832K�w��C3<`����`��V�WZ��:�O���g�W]���5��!��\3�-�W؁�	V�OV�S~���=�yEqlY��N����<���H#(C$�A U�S֛Z�2`���eo�p�YݳD��U4�ƴэ`�"��k������D����Ҥ�0�V �������$�Gw�7�5�xq���ˌm���V���|�"�����eǫؽ��#M���nR��x�8������a4���=�����s�����&)�(hk�|T�����xl�g�z�� �?��^�ws=y��먚g�P�v�ܕ=���:�[��d+��C�����":ӇT`Ǥ����,�W{b�a𜕕��� D��հ&l���ԅ+^w�
j.H��x�N���~u���͸q5t��K�rSRMǟ2��c`�֐T�xw@"�]�D<^I��K6��,���H	𜾥�<���H�X�Ϸ\�L%Ň��.�r.޹���}P��p��eƹe�.��b�t,$��|�ּ+�����6�n����b�3ؤe�P�v��.`��Ķr�W\��\�'�G��敪^�^����HB�,���ל@�x�2�_���0G�tVh�0��A���w�z
�^��0`��u1�R����>�8%�\H���� �_i�:�F��@��AD@�0�y�"�����vn�
����Eӳ�[Y+'�PA�u)�o���Zق����!2%�6{v�r ��l(�@�}��A[�B#wmw�j�=h;Ps�\doQ�>Cń�'j_�����\N�v��H4;����j��:��o�9B푈ʦuELlV�3�/��rc��.,��q��7���vT�S8�qF�g��v������ṓg?�"�����x�e��*H�g�6V����ǑF��<��4�F�|Q���hw���A�&Vu�ɀ%&.%7Wf�A���Õ㌐{z<��N���Fj�c�7�_{��~��3&��b�Z̘�Z��_'�m���YޚՌ��PN�Ǵ��i|�~6`�֌��u��]��5�A���?��V㰽�֌#>�y@���(�w�
��.)�F!�%GsF�a��6�Բt��cTz��ލT7�֎��¬6R7�T�KA��L=��m�U([|JG��jrN�p�E@?:D4Y�G� ��o}�{�{s;K@���T�є6��%JzA��X˲<R=;�)��#�		��`pi|�M$A1�$�_������ N��8��G�����=���-�5|��Ap0Ю0k�|��Pi��He6+�9[�k�^%ޜ|$˫l�2}^H�N���_�4F�g`8w�ƭ�[�b};�f`���$��+h�K%@RDi�[5Oidj�G͌u��p���� �C N��9���b��3pf#G���P��}���ȗ�d�r"����[�لr��|k�G�����e:�~p�"=��:h�u��N�v��y���7G���<Ru���!����a,�R��/oW��A~�ь���o7��p6��s�x�/��"e��p���<i��ť������A!���>�r�-�8T뛻�.��v����<��@�܉��<�%hX���Δ�'.tԺl����0�����ʝ�4qB�ށ��u�-=Z3�x���Ĩ�D٫jfv�<t�I�R<�۞\��nh5��$闘;qz��z����/V�	��#G�8��@_G��]�lb�=^0Z\ɸ�ʄ�C~��M������<�-n����%�}Z���"(3��@�*O���Rehf{�+GC#V"���:�(�:��X)ݎA�� �]�n���w�i��}�+���?�E��*��c�)|\m9M˫F���gNdf�V��2m���:�lf��� '\�dCf�;��iW �-��'*�:u��EZ�;������z;�i��K�K-i���aX5r~��b|�(����T�k>����X����(P����U�������*ח�9�c:@�^y,W�H���͙8q_j�<J��K�;� �bLF��	]�Kh)~j����w� k:�#�M�y���«��I��)�@��ֵ�O��UP��c�Ŗ@1'��$S�Gt�Se����K�g����%��M�6TX(&u�	#B�+V����Y:_S�����wg�S>ǎ�F�ȆqC?�tH$u�n��O����d��)���>t(&U��<�Y���x��8&�c+�n.Kbh�Qf�;l�#��3�w�n�*���m���K{䞲�֓�~�7���͢��T������ág.�?5��qa����GQ�2q�̣��.t�g��;��~��Y��/툯5LZM�!6����.�&�����Q<�&^i�HkQp\l��q�'�8��l.[�dQ�&am�DP`ޚM\؈��v)���6�OG�{&W ����d\��Y�K�B�8x$�����4U�m��9<�����a�\�вm>w�6N�{��s��o�;&�ɹ�u�	�u�3_�C��Q{��P��?}jF2dl���/��m?YV`��R�?���Bd�Ԕ��**���R��� �[m��'��؅#�q�&Ӝ|zU��'��˧+C�ʶ��S�)I��k��i6�ɪ6k��fLl'I���p	���9@	#����Q�|��Ef��%�53�Kq�tι�/^>fv���z��r-���@����4B2%E���8ɕox�����+`��MB	8�-l�^������{���yv�uWC� ��f`�1�@�"¤�ڌ�#@W�Q�Ƕ^c�Ć3�}���j ��zޫ]�P��pm�ii�,3$��g�*8�� <M6�:�5��>E�	'« ��!��p��8Ⱥc^xA=��|�QY#�qzm=��uu�����T0�"͚6h�_˫�����3'�s,m���� �0)e�z�C3�r[�M7�;B��\w5GWA�=2�Y������1�:O��)�$y��!�M�E"��1�����	q'-�Ϟ�w�O�H��1�O1;-!�[h����}2�y#�_tWo�g@1�]�2y6ǎǻ`���OR�ht�r~�c��>�9��d�sfA����	��$R�z \xW�u��ejn�
J�l�a-�wP��s�T_���"�k�QC�������t��G�lܐq)����5��Ac&A�c��~pJ(7V�̑ڥ`/H�V#o�>�@�Waq'O� FFYt琯:�V/x�K�1�P����0�֒�B��>l�'XdF���'��h%�G�t�Q�r����v�;���g�N���\6S�N�В6Zs'S���i�����-[f���`��B�Ϫ�z$3���)�:2���3a(�®���3��\v&5��D^�5Ԫ8?�Ȱy��P��I3��qfꊞ
�;������x��V̽� �7�����.v�w(�S�DP�s":<*.��T9�g�뙭[���u
���cm� w�J���F2����G����Q���X�S��E�XG&�V���Ȝ�|�R\;�q+�@�����I/��p}����S�|�	���9�B�w3�^�8� TC䞠X������}Ñ�P�K�C��Ѷ),��Ĭ��>�ޭ�TSK�o������g����_څki�~k�)���!��4����>����T��W�&���l�<a�".ho��vkxO>�ބ��Fl�*UKh�k#��&}��lo����R�r3
��5�Rn/Y{���j�y���n�9�%<f;�ͦCa��|�.�][}bO�ζ
�S
�HK��S��c���n�;/�)e@hN@(��n|x���z���G}�{�*�;M�U����Y ����JJ������
��&���#��J�u��[-�8�|��Y�Z�A�	�ՄNy��EU�B�'���F�VZ��o�������9P�Uh{a4��6/!�)a�����R7�~6�N9�<���Q2 �E�����"D�)V� �5+�79� ��j�}=������S��A0u�.�U���hh��wC�_�ySL����q-Q3Y{���IE�m����7ҥ���a��T��2L����_HmЀ,��+U���T��f��[�9DK�aFː3�ZtB��0��w������`4)��k�����:��Z�����zF��#Hte�#�Y�T�x]&��?�7��D9����[��V��Q�4�ܨǶ�б$��J�nڒ`��'q�ѫH�48���&�I��� �AQԁ��HȖ��O5Qi�Jtk~�[ε*ǽ1���D-�a�9�<I���>��Ù��}%�
�ժ((�L�M�7C7�z{7�'u�����R_n�-P|6ft{ U���'2Vy�2�R,��i�Zi�+#�s$��[��*�ٳ	�A¶�+�ϊ�
����A,�y!6J֪g���n����B1��b�B��౭���%��Wؑ)�> �I?�S�pP>,b�t[�c1�J�I7@��a�`�3���Jv��� 8Bf���5k��:?��!Ay0
��5D�i���4`�+(�r�G`?�("KW�(��'!�<,�,��ۣ��^��VG-r�~+|�gҖ�텆��8�3�
�l�a���bhVb���1�1ߋ��B.嬂es�'����1��
�>�U��.	�8Dx�'����J���$]��Z�O�_i�&5X{����x4�4<h�D��	h3�`{�aP�	�\��%����cm�2|a�~.�偛{�؅"ZJ��=�Y�< �}&��`�v1&���z(�A�*��Z�;�H��f�ءXtaIh������V�b�]ҿ\��k�R����p+4�P���wZ����?#l՝� �律,��ٷx�򹠤���݆�j<F����8��$o"O�=`So����c8��� E|&�'���Z���e�.����4�b�]t~�[5^K���[�{K�˙ls��@��d]���P��o��f�~�ǉڭ~d�HZ��ˍ�IS)~Q�҈eQ;�>W��b~���)9�q�^���SN��-�� Ӑ������YK��n�z3�q�=#ӷ�=��[��q��A�D����t�C1�D��E����)G�u!P��R+
j�}� <�볩4+m�����NE|a,�nf���9]�tD���X�� VC��g�\^�x*�� ���w�2����چQ]ݖ�����)�kc����I�@�5/C*��r��c��ǎ��Ġ]:����G;�'X �z��#~ƫ�2q�=�kT ��^W��x̝)]��#d5�}����vA��4)r����-�h���p���r�$�MoG����[ ��VTu=�����ρgKU���hZ!�A�\�����z�=%[��&0^��4$�S�fg��J����c�@�ޥ6����٣�C��#�tz!/x� !�H�o����ט{o���^}fJ��f���;�������o�N^�w�[a��lf��j`s�@��%�%q�4�����Z��5���g���Ӝ:�����<�H���Ժ�v!��5�?G���{��~Ǔ�������%���(�t�f�E�3-��+S��'�:��Գl��c�޿��FsHع��N1g������
a��j%,M�0�UO���;��K�
u4#;�}�6K�^�i�;���f+Á%;���~��� ~%d��y��7T1$��A��菲�/��j0�"�y�PS�@��$-F$�(ziCڰ��G+rB��5q�=�5(��`�L�Ղf8&��+����8}��p��Dp�WK [4RP�_�+w��/�q�#�,���E������l~�2#]=���}�Z��̘��5=�K��"�Oz�ŬU��w�>@�.�+x=K�@��8q�� |5V+�V��+d��3"�ڄ�1qk�E�7�I�=30>�{�]4��Z1�I���MY�BVh�X�l�J}�V8����ݢĂ��=(��/2��ɼ	���?<��o ����( �I1�J�B�ٕ��&�h}����I+��8}�a�s�{���8���P���]�����	1�2W{�h:�oڔu�5J�l�����)��_��$oG��J��oe����W�V\#q�s+�;WIe��-�L&p�kg�6C�
<Vv��EE�<���KT�Z~m�i�5�/�Ny{��v 9o��f��ڄ�I��j��%,�P2�+YA�0�9t�i�2����)tA���CLĪ!ڀz;R�gd��>���-Dݜ}%W���`� �d����z���V��>��0O2�eC��#z�
9����)�ٛ�J"�ra�������BX=�=���:B���'!�ٜ�.6�}[]�3ˢ??<��YorL,&-���|��k7m���G�u�a5P�JmYnE���HW�xb��Gl?1Ӆ����חB	l`wȎ�j�IY���0>�z����ˁ>��%TO�}3:Q6ۤjW�X�=�Fz3�g��і�/��5K�Vo�2-���C��yK��;f���_����!2p/y`�'��U�-ސ����xY�����k�{z��A�C�Ҋ�+m�����k���?+!\�ג��uUȽ�.���p���Ar{-�k�e�.�$����W4렱)l�u���"}bv�j��̬+c-T�l&�	ںI�M��[��&Z<Gx�(�s\�N�3�֯�2���Z�[�*�쾥ԩwp@y��(n����^-̠��a��t%�C�?����[I�9A�2U)�0�SÍ�Yxr�?f/�����%���J5��<�yqYq|���8�m0�#�ތ#�'6����v��p��^Kt�x����T��F�\Lh>�I�����:[;�'q0�?�o"�C�]Ӫ�t/�85��.X4��{����J��t
���RE�"�Tz�������QD���Jmb!�j42�l��dXv�0D�#]��`�"8���ŏJ�tJ �|{m;,_�����z?��f�}��lN��By�)Ylŕ���)��)@D���Z�Ta�"��8��4��8ճ������5MHA�d}���i����JF���;���"Z�2����8V3�UV 5�ī���nh�`����3�&��E*�*�w�͜X�)c�yK�0vyt_o��G���e�?��|!/�4%>C4z�������h���lX�&oK�Wa��E�j$��y���<�O{r�� uF�o�nJb�dm����z��0�
3,�	K���o �:�^�4��[chE�^��zY2w�,�{_}�.v��<�|h�l��f���%��/�<쌵Y�)����z��{0i��"ݔ���}IO�2~뜮nU{�����-?�-�H�&��X)�Պ��`����	̘���Y>1-Pfq�㼼Z	��-6�<>tǱ�� ���a�������,B*�[�מ�m�yX<���T�GM֞�OcH��l���"J}y�ܯT���T�哒�Q��[��M�-!R<gvU=��j������^�i����:�������\O~><�C����pS���˼�ey�9C�����?��t����+NÀl=l��,��1"�(h]i{�e�}�

B#R��-{���3G\�{��e
jͮO;��:+����6�)~���c@�cs��Td��3�u6���r�*
���RP���Zl�F�@�D�wnd���^cF�\�V%{�!sض�4�X�.Qɫ�O��ruL|-�(�Z�t�wgB-O��Qi1�] ƾֹ�E�ru���DZn�1�&3N��W����̈́��v��� }��cw-�[�4.����eAj��ַ-3�D����D"0�7�P��6��Rދ�s[c�#M�JMRw)b~�;'{U�{��g�¶=�QKҋ����E����U�^��� H8B.![yp[v'���3�Sn�ahL����� +A0�rx�=[�+f�k>�R}g)�4P�>7+k��V?��!�܎�:�MDv�D[�@��)lɸ�AT@i��ջ�S}i�M�v�T8���ng�r]���ד8�Ƈ�)t3&.nT+�,�ՒRZ%�d���Z���Q>	k�iT�@� �C3�Y�	yZ�i]����_
����l���nu���� ɊI��{�>�Ӂ��-����v=�xu����{3�{�̯���s2<S���+�M���K6�C�lxT(Ƌ����b�@�	��M�N4W��KX�����>8P]qD��m�L���i��C�`@��!�	ƚ�i�A��9\����0TQ�F���
�W��{Ŝҥ83�z���*\f���R5��)5Ex.ߋ��Mʝ-�2hM�]��
u4�Q��dw6��e�Y�f�ZF�J�?�B��)HG&n��O���`|���b�"$�p�L�|ku3y>���İU�Y{�ǽ�"�H�����n1\CLfń.'�;s��<�C&@#v{"�<dr����5�彝<��<8���n���̕+.�P�}�h��a>�"��r ��#5�E�84�!�N<,V��J�F&�x)nD��޿+�L�ܘq�i����g�ǡR��H������wG;�t)���K�S�jV�H�k`k�y ,5�\�4�7��.4id�u�4�К�5n���iu ���
�,)I6��n�!q��՚�O�;{��~Z�0�%C;�Qc3I:��^<�ӂ꿯
jFn�uе&��Q1�JT(eAՄצI��'���8	-���x+����ӆ��f9��V�Hzf�v���U�
U�|p����O�l3�Ɠn���65m�� ��u�dοUmZ>��@��G\�2�h�X�N_�0 ?���5"n�T�C�/��ܻ���U����/�˨d���J~'��vlȣ� )��L�2ft���%ǁ\N���}�����4	�F�=��=R��g�O�ڮ�I]�M�˥�$n�ҙ,����ɇA�B?Ne�ǭiM��{���+��\�G"]�8��+q���Lk�����!�9`���]���\�(��������N�X�;�Z����\���ң���_A:�.�h,bs�I)�}���8ʉ
aH���j% zS����&�=��^�O�S��9p������m�Ep�E�Bqȝ�d���傋���� ��Y��ԚY�?j$_n��I���A~�f x��Wڳ�wmE���f*@�����\Y֔1�#�ٚ�o��f���kv�����
�I+[�Ȉ#�-�lTM��M�J[ߦ34޳�, #���iNЋ
�aW�n�C���s�^t�+I�E6�0H����y���C\��˪z�H���4�o�҂ߥ������6����a��KoL�
�zn�O��o���O��<_�����|��@|�_����#�ŵ�v3�I����Uom���#�V֫�Ԯ05�`57+������ox��
4�{���},-�����nwJ�l��{���Ѹ5�d�����O�1�r����7i���PI��[)�l"ݢឥ8��dF�	�j�Ҽ�ƼL>6Q[���6�p���&�D���9���a�P�<5y���+d[��k���K�*{<�u�<4�����V�h-˻!���<TE|y������¬i!���}�pVM����d.��z�����Olt?�J=
9���:�,��o�j��n��4E�S	�u��C#)_"�,�(�;�g��~�XZ���W)$#��N5C2L5��o$�m�|��}���b���Ԑ�PP�=���[� �x�e~o&|��ͣ+�9g8t+���Rg��6t��_2C�t���}�a���z��K(V���QN@�q.�C��<ʊu#ݢ�l�a�#SŴ4�ֶ?�̝j�/W����ӕ�[�AԲ[�L1�
�+��ſ���-_�~�?�O��:8-�\��޷p�cS��<��7����W�����2͵ń��,�'��䑉L!ua��w�H���P�8/�}��To�!������
���a5Z��eI�>�w1��e��jh�IxR��_�N��ߧ�Gq�H��͟.��=?���$��DJц�@����l��F�~��6��Y5w�\� �M��+�l�9X�,��ov���,�i�">� qV�yޠ�wa�&� �J���<�EU:[���%��T������O|� G�5~��9���ty���ӤN�Z����T�sk�K�VKwE@�ɞ�������jG���
·�=w��Vf�$��'���~�03�c���`}������A�;�*F�eH%C�S��		��E�EW�a���Ö
\�L�^@�D��m����J{X����
�=VrN�n�P�2~���h�n���|>joj��ZO~�*ꛌ�1����}Y�f���f^�w��T{���~��_`���l�.�gc���W3�A	��}������d]j�e���xOt�@�
m�=�����g��x���.燫GX�Mr
����V�'s�E���(��w�֌����%ݼ�[�Gh�=�x�=*`�t�#�	�2a[���>�wT{�ڔ�5������X�H��ݐV�q��
�82�i,�۴�8^7�v�Ŧ��f8)�1���9�yf�˳}��"�V��B�|kO����} ��ۧ�8q�6NRgTF��
��n5� §�R�kgj�g��������o��}�w�-���/��\_���e]�^G$9����3Vx�.=Wk���[��R�� Ē�x��������8\adt��P/ŃN;U1bo�ěc�/��S#��	$�^KQ�ܩ����� �����'������f�E���LlH�I���U ��(�ȹ���P\���(�Ú�p.�?f4��-`�-�^V���W9��s6�!����2%-jM"�m�U�� O�18x'��ȶgH� �e� �>��)v���sb{Z���.>��qp���H�vc(8&ّ�"a�ڜc=u�M"�w������`V6�=r��˔���2��	���k X>UR�h�A�!��֌G���Z �G�
ΠL��9DTf..+��Zwd0�@���a|���,��ÿ���#x.Q��{����zӎ:�K� x�!Cc�gVS��`g��&���hN���S�/%,�q`gF4.�D�3v_�AE>q+0�!��Ia�,�����7�%u:;Jl�A9��h�4ݥ0&z���]<����}��w�!zr��0��P<v��C�oR�Ϗ�'�4��O�p	��x��l��q�g�����I)�r���zv����Ǯlg��b���R���[��\�l�~7��$G�3\{a����_�e���]V�T���
��E��#�x?��!�s���f��޲�4����b��6T�	d�	��NT/��	&�qO�@m��'�3O�xM���*c����pr(����b��؄v�;�i0<7v�,��
�Z��+Ss7���7��Q�I.E�8��KwՒID{T̯`���S@����鱁�)CɕǞ�/�]5�x���-��H<~��Y�?~�ŕ��f���-�ͤ�1n3�b�ϵ�6���2����LD�-)v��	�e�����(��@�%��32�M�e5J�U���鎯��5*�r9��MS(gp�v*:�b�<ٕ�j����rPU�w���AՐ� �N/���K�z=��H2�o�"p���R%�n�n3y�v-�	[�`��áUY	�^����-�k��k�A���G&#(3��n��ZoW6 ��V%? �� �qrѷ�?���`�=TZͿ� ~>DR644�>�l�CPJl�'�3G	5Y�:����УFP�����*  ����;��敫��ծ/�k�Z.���l<�J�$��L��Z�Aɵ�ts�.+>�  3T��$$��� -����T�2�zMeǳ��^��cL�N tP���HD�z��7i���2�Ft_�[D�K?O��27�q�*'��|b�l��tpN��o2�#;�"C�@ J�b�YEKG�I7�:��}�ͥz�є��6B�b��N�$�[Q�lc���b�D�ފ����]�΂M�^hZ��C�F��`9�����>�$�^xu�07v�@A{j
�F���b��_1���I�8V��V�L�Gc�D�lLA�ǜE��QA4c�#��A���0���䄀��o��ڈ隗��	���yАk{�k��(Z^,����c+g�w��m������TN��z�^RQo��iZ�H����Ki�1Nu���UI�a����')O۫{�(W ��h0�N��5f��Z�Δ�-`�Utr����1�����T�h
,�~W��b�J��0�zdC�w���]��r��T����	�����f?#"HZ���B|��z�B��F&��5%�9n����~Zs9��U@��G�a�B�!�t�|kC���kY�V%���rQv2��䮹�O�E%��9�f��	Go9¤ox[����1dN�0�W�]�eV���2A�p��V�g��0׺gC;��j�0"6hx���n�$�`�>!=���&�^�3�jfk�ag��5ෂi~�J���(\��㷊+U��ʑZщ>zz��X�ږ����>J�{Vv v[ �	��ݟ�&�4���O�\k�pF_M�o��He`���~�ʠ`�uF�������F�W s�c����\�r����(x� ����&ΰ3.�Ӕt�.L��Fh^j� ���T�!V(���Q����%�,3�_-�-�r�x)���Q.��5	�02�v�L�-��㶈Mcfx?\�-�L��C���*��{�`��Γ���L�0�+��S�-｡uu&�?�<R�e$�%�4�n~����|rSΘŴ��%|(<�������)��a)�n>{8�p
0��^��-��ްrG8�'�2�.Z����:ٻU��f^!�g4F�pZ�/\3����q~k�8s��|�^�;��� �rHŪ�,ш֟rr��t�m6X��(�/�N���oK���n[��X�t	4�:N��X�p
9�����5 ()"yi��*/W�E��/��LHu�U���2�T8% '�k��&rY����ӾЈv|�J�t� ^��=���� �bW��I�heIN�5ϝ���F�H�8w�ݶ2�F����J�`8�i�1�,[�x����E����_����ՠ"��)a�6�����"���t�Kv*�cޠMBK[��\k����-�����³S�y]Vm�d𬑧ә���>)���m�o�]���Y�X��N+Q��-�Z�s�8��C|��5�{ܩ��Lw��;|>�
_|�����l���L�LH��g4�\K؛tC����T���D�a�#P��I��^��L�������ǒK���DCy����N��+���m�1%8;�c���?��RP
�ͨhc�&M����X��_��r���a�G\��~�4?�����'�����W�B^�,�9*�<��ЍNO>n�J��U��"��^�zX����~�l�� \���Jr�!4�l�8��.;�@��hՃ�
Pz������>Ɏ�AB�L>�I޹C���s�w�]�J=�������?R%-bXuU��?�݆`��&i��ɠQxb�/%��PHyז����Km+�%��ArgW�80��Hr�p��|���9P�{|�`���"�E���g��AO^L筭5m�U&mȁ�Kw�EHm���V؈�%jk�B)��a����+�e���	Ò�A�FW�d-�L�0z����1�3���`��<�� ����h !(���X�#�w�SS�H��@q��f�ߥ��ߛ@V����0���j���O�?������Vf�f̀$E PK}��	�|��R�voա`�����k#g=ОEm��O�錃ǟQ��ĊJ!:h]x+�NX�5_"��w|��Hm�/Ы� �&�J6٣Zq�[Э{��0��Z�͍LP�"���/f8e:Ř��R�8;Y��#~���V-���&!c7���)���s�x`l��\pH��$В�z��V)���4�%��̽���Be��Wͨʁ(S{30�� L��zG�*�խJ-�^] hٓ�ۥY��o's���v���4��\���Gy��D�
��®�'$5i����yغ���YK�U3������~�hpe��u����Þi��
o��:��Q��|v��x��$'����\V�h~�:{��N��/9ͬf���!�ɏ���X.J��?^�Ltzd� �:P��N�����dcx���R�h������g����+f+��.� 5Y�k�2� 4 ���������qg/����!�K%4���� �����/<IV��36��m�;��^�8�$G���],���੨LG��zb�o� �8�1��@��U�/i�#)�+^��-�"i�� �Y����m�,&�}�&������5֌v$au�A�Y��1�\�!g�iC���:�&wv�I����]93��o�d���7��NF`���6&�.[����2a�����* w0z�Sh��h�5v]��@l���8z��̝�����c)�I�G�]%ʜ�3߱�]+�P���WG*� ꣭�r������m�:�����X�!Ұ�Be_�,���ֶ�bI3��� N+v�J�l����,a4;��)/�g�R�6�4��H�͸��7b�a���t1�l0�\�M˞��p|��x��G��L�da���#yX�~�Z*��!��!�,���{B�4��9!���S�	��b��t�Rݧ�	��KY�=��E�"ef���p1%#�0��)C�f��$k��%��a�L�����2���W%�LA��(F�|�cd��l�z���_���{�	�Q���h~�BX�Y����a�↢���P���~���+�,f�"Ϻo* f�D�x��o<���F�����b/jk�ft@##u�:�o�KD'��ףҶ`-}W�Ij����*���&V�B�XX�C���T��L��>A�zД�@��/��w N�_ӷ��yjP㨪j��
�.=슛jg� #��oT�6�Iw���VN;1��v�:9"@�H��3�$N���Sf�0��B�,�?T�{?�H�r�Kc��	��Ǹuڌuٸ�%����̐H��P�0�P�zP��Q�!Bwu�Yu�`W�qTW���&S������ c+c�~)PE|I�蛭���m���3�-;�u�7b�R�� ��x8Y�Ђ���B��%�2��&���mI�a_RQʚ`&&��Og���<j��Q����6o{EȰ�y�D|����IvU�s�f��
�CĆ���fDY���S>�i��3���\Zx�z�V���G��[f�"�"" �%�X�X^��8E�I�X�y �T��no?��:�t���r�-E�0WQǕ�&w�,��-��U,MB�E�vꗦVz1��/� ��4��-�b5�����L\��T�� p&�RpZ��`}���6�5I ZU�B6�G����K/$.�ک+�Ʌ\ç�"�i}�(�A?Oy��A`e��Te��6�<B/���u@ؠ�r6����@���j�����P�|�u��ƞ����n��47���yo�D�9�9���:��9|�_�ȥBK�t0yLc� l;lՑ�)��o��_f�f��e�
W�����>�rݶe�s�=c؎�hEX�V�e��2p���v��3l�o�ͥPS��s�=
&��g�5�P:��Q�to�ў��u�9��l��O;������J��M*{|�ǈ�U�<���
�3���f`�����E
x�>� �iAΎ�Z�Αsv������7#�l������5��\��� o��ѫ���R�2�5�q� ��v��5Xϯ�;d���и"į���2Ό%$"l.D
Q����qGMDV@e:��9Qc�v�f09�l���B5�<v1�:@�!��{R�wCwJ"*��5����g8�B��%$;������$8���.(�RY��j%[��*y]g�@�Q���CA"�M���:������2���)4	�Do�K�u�`*g2�<D�<����iXZ�׷�e��HU��O�iv�?%ֹ��umԺ��" �=[-z9N8�OL��oh�������.��/4n#1��j|��O��Y�hi@�~k�^\IR���|��	�5���#ܚ"�m�k�cCܥ��]�M��s�_�3H��
+���|��\O%B��f�
J���()�	6�v�ώ��-�50������LX��.ܚl�!��`:��t���,4�ŹxV	ЍV�� HG"Y�W�gk5S{R)�w�m��0G�3Lz��
�K(�x*Y�X��5sh*w\[T�l�N�Ie�mw2NM6J*���ǵ.�%YJF�iT����8���	`;�JK���:���L�Ks9�[|�����Hv�H�
/qW"��fa5d��:�&wB��2�8�/nj���
Sq
=�wڨM>���U9�I��nn6�W��+������i�\� �i/��n���XKSN\=d6�y��Wr�Di�J��]�T� ]�@�Vc�m�ދ�#�ӓu@�n�:�Z��E�RC�Lm��8�+nhE\ o�����Ia|�!I�=5�8��Ei��9c�:#B�M
�Meh@H�gx�̍�2,ko+S�~����:$x�\1��#��~�N(skW�5I��$ĮB��hߒ���}{�ͷEX<z=ߝ��`� 	�I9���Ӛ�<��T�)�
��Ԛc�S�:x�ե)�$�d:d�Ͳo�!^6)�P��2���]��\k��)v��?a�r<�^�l֋���k8^2��:��j��`��rƺ��Jo�qrb��D9��I&��Qiܯ�m���3C���^�-!����m��=F��R=�Z�OVTڵ}y1I��A���`��\с��jVY�!H������C9^ b����J1Lb��Y�.��`a1A��q�2f��Y?��V-eugO:}�^Fu�l�^�(�ڴeBvNf�v'��38�M��������x��v���y��ïf�igo�B�'��¶���.ωYj��(�+� B�%�1����$l�O�����cU�~�ro�@<yn��B����&��X�P�!����c��m����.�2����L%%W̘��ԡRcg�j��y{9�$��n��W B�L��&�V:n����v]o���=ǜ�4 �1��ZE��5,I`Ж�X'S[���"���Y�;3j����:W1L�1Cˁ_�4�P��ټ?M��B3pu`�t�L�=r��XeX���*�Y�* �`���=����ލ���o�_�����2�-ȆPg��^��������?� �0$ѬT�W�����Dj��	JW0��a>H$.����J��<�C��%�I���t8�6<�9��������C}n�v��R��z�F4%	�#��,b}�]꽪��G��X\j �){�Hd,�A�#3��
�a8�H6��/C����";�wL[����2���y��o@=`�op�ȱҞ��!'� � �|B��S�Y���B��Wa�5�1��0g�?�pD}̪5D�.��L�)$D���&їz��*R����7�4��ʎ�O��T�߷HQ�Hl�$K0�e~��*URKE�˻m���8�(4�˵=֛�Tx���z.Kd�.J��
P���D�|�n�Ɍ���xq��;d#o�Dn��a)�vw3�?���5�5U���^�ޮvƈ;İzʓ�!}���`�e����|:���UOzۍ�W�^īN:#�2.+���X���LX[�ӈ��Z�}�"��N���.Ƽ54����R��@�3e`u���D���e��2���m��2��f��O���:�	=~\��uӲq�RU59����cB�V-�d�[��R��i��\���H���SI� ��cE�9����&�b�Kj�%k�
-P��=��|S=��X�ĕ<5js��UQ[:���5�~p��@���i��j�w��`A��l��wػ�)/�m]�U��wDJ��@��ə�x:E�^^Aq�t�g��O��U�.B���N2?u�]ޑ�A���d*A�3�h= X�/;���1ep����Bh�u&'[��,���rG/�L���<k����6�:b��`�tE��˥��"_�UA��0b�Nk&il��o�VX�3��������W�F��RV�c7�(;��l��@�qb���X=�[O�f�T����nЈ�o�M{�����Z���9W�l(��ݢƟ7��Ճ��]���f��~7E݃3dj%�DJ�e$�P�����L��2�>�nBSc(|ϯyD�[�	����<b%q(A�P��e�^��r�mcDr s*YIn͓�+�|YEW(Rߪ@/�O�qra�u�A7�Pf�uC8�ńL�������o���3"ƃX*T0������xG�G��'q)X�W�(1_���2�=�r9.g<�fW��&o�8��J'�X&N����p����ܺj*rL�N;5@�ה_�����W�b��j3kAUaa��S��Y�mA�b I8q`8�Z��f��9�W�7<��D��S���O<�r@Cl�i�F���-2U��c����^���!�����eMK��A�����3�H�P\/�}�]��*��Ux��0u�}�^@-�b=Ir��O�n�Ǳ� ȵߒ�Z�҇?kb@���}�{��ڗ�Q����W3J�#���)z拈��)�C��U���I�zs�p����iCL���)�p����h'
Y���r���q�U�E��-;|��8�N�!��6�.+��ˍ٩� ��X���c�[����XQ$_�Ŏ(���ݟ�H��Jߛ���J����m����ܤw����S�֌���c����6TN���n���R�~��ź�VM�~>jI>7��]p�=�$?1?q� ���Ba�fn
�?�s�⽚hm"Et��S#�-b�`�-��_l��P�m���7��\3n>��_�ci�j�k0�ܨX���"e�a&vKó\{�½*MxP/�ɘR��Q�'kv9�6c磟���}��'�>] у������M��J� :��@����E�*��"����e �c�"�<O�r#�eC@�L�C�(	M���*4��b�nE��%�U��ŉ66����S�W-\����A׽YOF	#rc.�0\ ,��i�ҧ��e�B�N�0:�����GM:�]�p HQU�sV[)D�4V��Du� �����>O�R�h�����uw`� $ �V�T�������� ]ۀ����:�
��ܷ>�P����P� '�����BR��)��Y����C^X�_y���5��S�ʀ�eP^[ͯ:=LT�uK����JmD=OT�1��w�ƸH���+(RO
�S p~R�����+��p�0����(H'�M��x@{��dʳ�[V�l���0�g:U�eX���R��]�I���ְ�a��,bN��e�)�d��Q�0����\"�q��0�ƬMk(�����?�	v;,tJ�Wf8����<���5���b���0)s�Y/��{,p��mD�idaJR�$�|��[^�{����ű�6�^�̻<�F"�AP�� �_+
g�by�m�(��<ex��A,�5���n�����_���$|���*+����ac����c~y���i=�Fܚ�d�6�d�+�cN+�OUk)�~I�6������&��������\d��b��?�3V��ߋ�w���E.,޳��b�����W-�!/�!̱��</�y�P�n���D����~Җ3Ր"5��d��+ղp���E��,��+��y������E� 0�Z����q��_�Љ����卵$"�%�lf`�ɱG(��8��q��$�`���^9o~_׃����HY)ҡ���%*����^���'�4jv~���3�k^�r{�vh<�ӸjN�t���:�$���:��8���r�=t*TO�X6٪�4a�������~��Cd�����L��%Y(IĬk�gX���<%�.K�@��ªQ(@�d��IH|�5B$���]a	 � 示��0��ϟ� �j���]����V�_=���Dq���X���# ���~����֋��
絽�x��C�u��q_Jw:��)-��e>�B@O!F�Τ�u�zqeM�:a#u�r�j�� ���k���|CK�թ���Rs�j(�X`�ȯT	
�o�G�.S���-�r&�3�VA�B-���R�9?���]�6�,�oynC&�t+���y J@���G�u��v�Ȭ����IQ�$��Kb3d|W �N/�Z֑��mfi%[b��&B���2#C�)$z��&�lyA�,?���ӿn2$7�:��Y�4��ߕ`9�!�a璀hh-��<�z��i��yN%t)Rk1��r�|�P��G�2�\��1�?��H�6��V�4��`��ԍ�� ��>�'_��dK+@�Ei��H�!u��1H���p�;��I���A3�;�0Z*Ҫ�Db�S�g<ᕫ�����dx�QX�j�K=Js�D��St@#5�ap�e��ψ\s(�W�͢-q��$b%�����c�'އ*�W�cR�ڽ�i�-{�7�����E��3��s�^��r���͹~z)��3h�j�D��ZH9WW��P&)���P��n�9��g�\>���Z���z�۱YC�����7��l��uh�U�\�U��%T�.4Ȝ�W1�kl���3�ǰ���v}�.p����8��d>6�W=؃��.��^��A�JM׉��I���P���ܳ�'���t��*�+Qa9#m����%;[d���c��}������������ݙ-X�.L���~�V�W����;��n.�?r%MĂ�Y��.�]�$�Q͌%  #w�D�cP�u����3��L����yz��LԺ"�\_��`!�7/U��T���.W�;��#N�+.��c�fḾ!|ٴ��%Z���S���;Q5���
��~�d{D��.��ct0��f��L޾�xd��jN|߈�s��%�q���ѹ}Fl��b�o)����3�P�V��'��"I^ã� �ϻN�a���|/�joK�w��3ΗTi�C����:�V�-h�.�p��4{Z����U(��a i%����]<��'J�)��ȦO5i��7N����D�I��ۋD|�,_�x�ʕ���L���޾|���E�3$�:�3s��EB@p ז��d9�4MUS�V�>�(�Bv����@�ۧ���g��P(��[C5�6T��a���q68��D��r�� 9��MZ�̛"��"���G����p����H�Uz�Ԙk�#�R��іT����[.ޗ�fU�A	�/�����T����*|=@YrN������s);��\�L���	�d� 1S�3)����&7�IO9��uI}���q���B-���SD(0 � �D���IPu�5Y~��kS���e"g,V�QY�t��ճ�Fd+�q~<�l�C����D�P;e\I{i{�#�C$�W�l��La�ua�3��o�'�ؾ��\�.yxiP����殹Hh��4I?d�a�ik<x��l�f+q�0�e�$o��aؾSO�v�&���]!���rmb8r}���T��z��..�%��vE��$���G�j������c���[�m����a�D֯D:�x��jz1����h�uռ�^%�;zB|�6j]M�*n�eNhՓ��=�3{BG���&�I)Q���h��ƛ�;ǘ1 n�?W���Q\l_����& 6�i�֛L���J0�_�@����yg��k]�Y�f!s��OJ79��m�齠�n�l/R"�8�kB��4�݌�˺L��)����Go��ʤ����aL��z���9i��SU:�T�'��<�L��C&Xa}�tL�&q?h��I6��l�3@��i���&}��/���po���D�h�fx� m���>�#�y�OfL_��<��a����Fd�m6���Gqv#*j��c���$t����a�xķ��^�FM�X�f�)��z�٨��*4��`O��b"\ ��Z�["�� ���z��9}�
T�J�&�o���jBp ���q�kT�zH���F�~�Nu���g���	��4��x����[�c�FO�c툼С��2E��n=�vDK��>���.�kΊvH�-��܌3cֽ7��4Ǜ>����s����p���wv���"xD��#2���%�X�i�b���Ü�z5|`+#�>��_����0��.�}�Nޓ��9O\���� uVXt�dNݏc��ϧ����
�+�0���`p���a�3�s��r�䩬�ܼ��Q��3��]I�{6ߕL��d�g�\��;g*��Sڭ���;o�Pw�m���$K�hco*��h}��V�bʙBs�8��@dx��c��+C;G�3�c�ãU�{�Q#��+�^����ԻcI�6�1+"��8���L�}�mB���W�OWh��ZM�N��<�x��P�9���#sv�-�ږ���S�Q�-23�֓�x�d:څv�  �9!�x�Rh���W[�v0�Z%�Y�(`�e�e�ʬ��b����[�-�����4hG�� .���MK���B���M{K��@?�>Ȅ,�Ҁ�B8%�
}s;#V�0�cvt�^�:SهՅJ9���q��A���%]��OW���L�v8?zb=*�.(�ʷ�����r�r�=*�>��'��@�{&�ԠXӯ�~��(�g��k�|q����	���|9�\��}y�)SZ�Bz��=��PI�يS<�oN�Z�=��O �GM�	#�����i�
�]�Wmq�_Iy���ͅ���f��N�[�y����$� J��9B���a<{�I�Y�Z	9?��e��s��՘��W���ӫ�t1�+![����s_R�T�e;�bX%x�b;/�^�xC��&5J��`�'	��&�~��z�]aF+�BQVYϑ9�;l���W���!^5x6��ߐE��鞉��6�{Y;��1�9�?���$����*�r�8~�1Gi�b�d�
l��H�`6�������8;!�B5�&v-�I�#`Y�9�vzv�^��p�A����� ��V��� !��F����{�W}�5�An�=��p�
��~����#Z�k߅�p������Ա]����ل���(�\F����C�"b��"I���pIF��=6ѐ��20��<i����Z�h�.$_�	ǆP^��)�a��N�{)�x�϶�F'����	`���֔�^� �U@���E�{����6A�H��v'^1�'ik����"u�p�a%��XPfy¶�_����Idt&crݦA춋�����l�,�y�bo��kU%�4��e�?���`�c��*}=���d��2����̒kL�|��>]b&�D�gF�@�N�??BZ�"y� �3���޻t��x������H[Y�%h��I�0G*{��M�h:��tu����c����㨸�-���K�gz0�� �T~�:H�ve��W��?-�y�S�P�}$ଣ�iwT�V��w �A �2�`Tl�c��P�Dڊ-��ԏ�	��^aZf�z&{+]����g�	��TAP�6�H�+ �l|�Y.�T,$|R�[1>�zTw��֬��^��w�fLl��/�!^�������+��v��d�賜*�����+���ko�c�_t���Eh/i����ש/	U�'`<J��r�L˟ͫ�:�roP�FD>���_�SM��4�P�z���U����/�!�7�<���_W˩�ӆ|�Bc3g"�(9?��zvYK��$kyM�~ӹ�Wk��܀q�gX
���w���a��]�7��Y8�P�H�'�X�I o�ϫh��|�^��a�5՚��8�]���r0�y�צ媙�.bң�F6����}�X�x��6���C����+�%�P��0��E���������2Yl��<4�<�)�e-s^��\��ډ0�S���V�&|F6K����}晇����B �hG���a^F���:���#�Z!�,ɔڔ��*b,�\,�p�IsTu_�d�@�tK�w�/s�A;�����o82��������5h���!O���N�1z�(�cH @����X��>@�W���B�s�U{�p �4Mc/jqq�e�nTi��fʺz�Ȇo%[�̀^`��9z��!w�GZ9)�{�fy��-z,�T�F����p��a�De
���E�����j1`P�[���2z�3Ƅk��zn�����L �3�)�遵�9�}g�-k�!�3.��j�*���EZoo���X�/�[�4�S_u7�#�� 8K2=�$ �w�p���$X?�	*E2?IDt�g�ǚ�3%7
��1-eo �c�R!?����'p8Y�O3�#�=҇���%���{i�Px�V��  N����dt��q�`�N�!\�{
K�~Q������U	�2 ڄe¤�����ȵ�;�;R�]j�A,��(�� n��k�T��OL�s�(��.�'Dr�le�z̶b_C�4�BVR%�5;AE%g����{D�vA�T�۱�]#�e�ڶ����];�I���P<M��H4���/�?����;���뎃�"~5�*��6�_H. K�JI��7bù�1!�5Eix�'����-5�^��]�a�� ���1M:̯4��W9f���]K 0|I޺'�Їft�(�s1��S ډ�u���I٦��<#�-�~ZwB�E��+�������av5(�:`��NH�~r_�`)������©�.�z�M��g��^��sm[��1��ig��,*�BV�$dIm���4�`��'*3�ʸy�/���藜�"KB�HS������>��A�Cy��i�E���{�t�U�Mce�c�3 Յ�9iމ"�������1 z�qߦtws�l� B�j�މ3E���g��
�K�� NI9��CF*�勸�30Οy.$���+`��F�;���^���L���U�t�˴;�zb}[
$U�Fv���`��°���� r��xq4�v��y�73��ӏ�l�\�"'����C�#)�éS���<�{�"NI@��A���6CVV*^�g�����8���vIr�(i>��xu�%���3��MM���t�*��j=�eq	��p�z3�/��&��څ�xf�X֬-�~�&���f`U�s��a70�� �%��}�fO
>p�r��~� @3� A���|���J6��=�M-�£U��OCS��U���ʽ�}�B�J�+.��������e�6�H���+~��r3�`})�0�g܍���NX?�������.�s�����#ٿ�AQ���a1���c�mr�gq�\�殂mI�sFawk}��0jL7�Q'�5�d��E��ƭ��z��
��x}��=�K7!I7T��N%������[�|ɿ�j��cv��V�f!��:�}�Nk�iEא���3�˺����-�3O�X�ǫ@Z�Q����֏GÎ��%MD��Y �������JP�9�����l�4Ԅ���<v�Ҫ���%u?�h�V�:���l�ڠ�o�����2x5�c}ů@B3y� ���!�� |���w=�� 5� ,�R ��g�>�1�'�m$��n�_;
 ĔȄ��y������ة3Z<&=A��WR��'��$�ᗂ��3�Ҁ;~U�3X��R��t;gc����^K�2�_z�����Gn�dִl�� ���ڒ�IFt��v����Ō=��qk
ѱ }��p.q�qW�q��;r���;&P�Od��L��*3ZZS��	���#O�֗�ט�1��q���y���e^?|1��,M�Ts��PQ�FȽ�������' Qi}�Ԇ%^�@�wt��!�}�m6H��d���4� ��9b�+yl��*d��:�м -D	?}Ѵ���	��`��� ��Z<�	rN�W��b˄��m������35w8�&��$PUh��Ao�Lݰ�战(�g����("u"6V�)EoD#Ǵd��ry�Ei飆��\���t�����À(d�xI6\���!H���N�wR����S�&��
Q6?q��A��?yhe��
y��h(oV�O1�Z�8O��F�Xn2&>������,C��7����l~�ф�>fLnz�ۥô$�$
$Xߕ�VmY�AL���[��0L�ֽ8Xb�6�������4�Jz�wlg�#?��	Mܫ��M Aǆ�5��� ��"��]i���m?:����9���m�Mk,%��$�t��!�L���q��K=�W5�c���.#i������K5���n����:� �/����V%zNj�}��s?t��ܣ2zv�AW�g�bۏ�M)+�J���b���)@I�e�M����9D� �LW0�`��Z����+�0��Ւ[K����x}�t���Q�%�"F���'m#�I���͙��ZZ��t��<S�J �;b�����Sm-��/���T��v����nj�	ɸ^W������0����sh�Ά�����#��nj�Q�d�X@_��`�����!<0N��<�4��)�E�#|����cOAvZ���(�ƖOe����Yݪ)��$�[.�����j�Ę-�B�r�v�/[����8�BS:_L\�T�j�#$`�xTî.9���7����:ㄼ�� ���k����t8�ȸ���4[�Ȏ��qh��Ь�E��<��N�@]?��/Q��\|��:�W'�eH�l�O��dL��n��fM
�B]�U7~L��_:d�NWP�gg(�����^�`�'��n��OU��	,����3]�aUv�����%.�x=�s���q�/�b�ݝ��z`��n_,rO���٫�]���}7��8UW��HT�����,gE����ݍ���!�{N6R9?@T^l#%54z>��ɾǔ�dK����T}�s~��$������v�*p-\I�_I]+�۳�"l{=r�Jl�����S��-�
v�
���k�D!)b�ڟ�^<��NLg��?}ǰ�Yb'�Lk߭��Mk�D�T��+��pȧ��;�J�6'O��6��d����2┨:��-�(�3��j����sju嶿sF���_)�</}Ҿgf���yS�T�"�A==����f�x�B9�6�]�gz�ѪI�N;��l��%�v��7C<2WU�.�g��Z��D��W4�3��8�uG~�	��1�v\�A��2�5��S��k襲4�D�[���z:����N �Q�v���������e����q�
��^�[�"P���1�}��7�il��,�l(�Np4Y��l �4(
@����,�6wɭ#�92H��\��cS?��8q���,�2ew�V��G/�a/��r�]IՀ�j�t}�I��%ݧ�VhX[?���|�h�̕"�)%E�;-��&�	���MX�^�燿�U�Fo�Zh����UUƓǟ��_r{�2g��� r�N=m�f�Ɲ��Z��J)i��O�G:���v~H�!rR����'�QK�[�(��6�x���K��$�zrŧ��m)�&??���hz:�jh�&�r����D�*q�s�r��R��:U�#�'�T�5GÃf�(mb��ԶU�<32�|�f���8ܣ�V��0 7��n��I;��WS�?;�e�b��I(N>b���f|ƕ��,�eI�K�����Q���(V�Uefܮ�h��2y^�N>�;���;�ʚ��~��;#~$�jN���̿�0��`� �y������)?�U���iJ�z*���e�č5g2�~��}Cg��Z���\3�*��D`���@ ���M��ͦa�-��v�*��V��H�2݇��^Z)�v��ͳ���ZZ\������M~�+[ڈh1�3FcYyo�X�h��A\� �G�G4{5�_\�#�����y:x�s���0\�  Xs���+�L���������o����@�Ox*�t��g+j��f�ei;�y:�OS���f�Q�����&q���c�p��)]�R(�SR�7_緇av�����#BvU'�;IQb����Pfo�mO�W������}�kg(��YP/��F�P�ʞ0#��?�C��.��6L0$�����~�0Y{P��kW��
�i���I�/��n�� q����=:S����}%^YHL`ذ&L6y�/��燈}h���D��L�#̘rM�������}�J�"Vk����z|1M��W���[��M��R!��k�5��-��9���-8�*0H8x�>ymQ�⑁dR��J�]}3�!��H� /k�POe0#=zū鐉9Ą S�{�l�bގ�ڊ����y5�,NCW
����؋#%,����İ"�JI���� ��v���9D�IT'EB_?=`Ȃ8����
�� H�%�g�m���TM��k���vܩ�|����P�ڊ�I1���"���[��_7���|&�H��r�2��>I�w_?��es��m����$f[_�dXIR���ތ��|�a?���R��3E���	
.?�jo�L^d\�|����h��mp���^E��u��9�hP����! ت8
��x we��^9����|���c�e�m)'a�#�]�+��x���\(��� yt��HQ��L�m�Cz�3��%ԕ�lC䋼����Z�*�E����A������z��)cb7��ZKmȃ�c	�Y����9�6��/�r��������b��ˉ�����<�z0�I�`�a)�?
��x�+l�C�!)�M- ��g�ݎi!'��/"�I��&���ދ" ō�ʓZV���������?(�̻�[aŴ���2{�p�;�Π���4N�5�¡���bZ$��/޳�;�[�a�s��5�j~�3��FNީ8�M94�+@��Q����X\�x]���"_}��	�4���i�H[�:]/qKo���6˵1wk>����2��@j�����[�����h�e�q����r�w-���8�,���/9~ p2�8Z|V��d'|�ԑ�Ǽ#��pI���i�i��b[����:����������X���M�HiS�I�l������5]d$`;7"�5����G%<�:��Y��4�_�Q���	���|�)��Ȕ�XTS��[���7����8���_T�P����!��'>|;�8�t�lb�_k������1	J�1�a"
@T�f��S�c������I���9L�F6umj�2`b7
�ޣ�Z�Ǉ!�>�_)J֕�Lq���q�/d���n;���\ژ�H鰅-��g0F�}a 6ɸ�����q���J��Tp~�{�2�e��(�d�zއN{��A�}_�O�ut��N�� m~aˋK1�eA�	.�����7A��ŧ\1�
c0�|���:1�[�Flr�Ю{@8U}� =�bK2�{�J�������gL�<
�{��$;y!����'-�>���1ɕ���wp��S:����o�h��'�=�e�4���Q����ˉٵ��J����C��%^�Ӡ���(���(��)�7�,��#T��M|������6�C35�c+Ye��s����B7H3�˟8�C��K��y,� �8#^���8G� J��l6!�P���D�9#4�	%�?��tn:z���Mԟy�k�� �*��W,�!��Τ�e-1a/^5�����{J�2`�Q���kP�j�}�$��Fq>����t������Iț釚����ܫ�Ym���@.i<�n�(�=�D��bX�������}N%ٜ����2�'>�����x(.:�3���aF� z�yQ�N�M�DA-�}���n�|'I�h��2���q\��U��@��j���@]� +y����`��W�T5�G:e�� ]���Jˋ.�vKA�L�^��.��
v��XD��_SP�5bz�B���`���5]w$s�8TU�Yo���ڢ���`Z����C�� �%|��d��8��q���y�Ka15��N4�Wrn�5��~� =Htsh���ɼa�/y���F�½
o/�� E��U�3(��[/����,���oբj��&���<5�B)p�۫�eA�=��3Vn����lN���_	�M�HB.�O�2����"^��=��Ęox��Z�?�2������)x�X
7ެᄵ=?��Ѕ^N�=S8H�M�dE�hyZ�X�D氲+��sn'`�S�D^��]�����Z��k�Sb�!�O4:r�W4�˚�bQv����P�t���b��M黂�i�GZ*����r�6��O���%��~�|�"-�h�'!��ItCy��y��ڜCS%Q�1�1a6��qX*�	�2eWW�rooGX:	2��G�}���z�Tl�5x��^������v�����=��������Z]�5�(������`�Ĭf��
f�8�@!��F�����Y���G��!o�-<���^uP� �*����>.���\�z���/"��T\*_}�<@�24y��̉�  �3�s���;�L��:�W2��Ԉ��v�l��W̅���@�P?��r��]��p�C���7T 8��J	 �N��4C����lE���D�
(�&��?�������P��W�7�ej�{������ d�90C{��e#I%��n�l�A՘�3���4��m�yh����c悬#'��Kr��Oǉ21};8�&��I�`�e����Jʶ�,Kɯ���P�<W������&��Z�*��v�>�K��}�k�����(@�s��KZ_���m�E��d�#���ٛ�ct�׮�֑�y�T���x�'s�keT�E���Q�?���yi�
��5�v���������XU6��� �I.|(*/;�<�a��q^�mI��do}&���l�H�mU1�O:�$^:I ,���i���w�sD����j]j)��x��@��u�Q��|�0��?��F�e�)�t_�sW��*Q���+��=�D:�P5�����^��累NnBY�k�:x�O�V��-~m�rEK ��` �h;h��Y������+��F����RE}�['����e��c���H܄�0?ę8�I��$Y~�'��xŐ4���ԩ(/���J�%�����k��n=b���Mw
��P�CICE�e��*���xR�@�5Q�ˀ)�l��|�6�n���B��r�Վ鸸�~����98���Ζ@,�{��hhk�4�*��3�j<�NXy?}�Y���m�u��5R�4.��I��PO"w��F~��pG���>��<�P����D*t�C��zC�h�t(ҳA�Ԟؚ� $k��%�ME�k�!{�s�
z������$�~��� �ߢb��@��O!� �9p�UC�knI9$2��5�월�c0��GCDL"�N}H厠ti�fҹ��i�޲1�|	��-̛+��Xsj��ðU��iU��j�)Qh���[�%����<����e�X�$.���O!)F~md��Jȴ3�n��ו+�l����%�D�F �:3���
ķ�E������d�tT�ްz���L"�6� ?�p?�M�-�p��g"�C0�;�v�L�9U�=.'ߩ�R���U��������G�۱�ϸt3��ğ��f�bo{|Q�?��:T�O8c� ��?4Ty�Ń����V
�c���f�D���eI�ۘL>eT��6gV��.�'�X)\�C�����]�7��}�����r�'�:&md��#��s��)�z�a�� Vn��iYrgh�<�A&�'�{}�d�gk�/�՚��ЉbGԱ�?ͻ�������cQ\ �"3d
vc�NMY�﬎�7��G�m�����x|@��e��9f��^3V�0�Epk[��vl��iN���ݤ#=đd�0+����\��w7]��y�&ڳ���;2:�b��2�a�%q���V�|P���$aMH�����F��h0�uN�q
�Ʈ�`����ƺy0c	!�����O>�C��2�����
����ݓn��+yx��'\�*����yA�-0��ny7��.q�,:]��P1�	� �:<�4J'��X��N�rv�h�YTt�l]�N��9k�y�`n���%��M�[TN���@�'N|)��f��J^[��K�;q�*:W�;����;LJ>�g=�$�+�'��"�F��51+\�&���.�2M������c�$6\���:v"5ަG:��d`Z���?�v7Ө�����+LT|�l:��g�(8�˳�v'���%q~/+�R�"D�ɴ)��ޙ���S}��3���Qɛ?�.j���/�@}j��̿�S3��A���Z@��!*()�����Zi3�EikXp�_�{��Hȣㄬ�"oc�Bq�߄��Ә`|�+��j�� \3�(S���<�:̡
��O�c�EB�F_h�"� "|y�/�`b7P���`�,����*�-�@�9��k{�.Yñ�˪�J%>Ș|������N�G�y�:X���/�"J뽵RL�͟��>�b�v�3b�-����F��o\@����J�>eZ�U;�$+(m�W�z�8��)o݉��Sb�7�5]��SL��P�J
(�4��X>ȵ9�Sh����M(�-b9'q����������I��QWB��<����k�%�R(|ր8Y���p:ɐk7l�W�s���Qƥ���Ի��l/����dp��	���P��AW�X$D����mw��*�J��)��·]��v��Y��
5�%��k��Qq��n������F��X��"�\�aS&�_[*y�D���#�'�rD��s!`	���fm�2>�Ȧ�4p���]~ I���0��m��G�9�-���>�n��id=�`�p�x;Z�q��JS���sK���(^�dTwU_2����k��i�0t¶�Ǯ�HT<��Iu�O�!ĕ��^��H">�Ԅ�!�W�$ߐS�c�Yf5xp���z� �9��J�̚��+AUb16�Nʐ"�t�X�	�@��6����f"��C�N�	���&������C��_��G�)�^(s���F,dJ���h<��x���&�m���bA��n\'�����u9���'������V�,"o11��#������;���4h�����E�g#2_������஢��{��,�jE�$�˅���=�|mmWȐS�IY���==Q����{lI��hvx�	}"J*�h|���S��]+��'Kn�0��{�������	6�c{W�<���3!Ks-�Db�XY^w؀�/�����
����b��y(R0~4V��DC2*&Zp���s�Xp~ n�� ��>\�4vjA�cc��c��ܷ��ly;^\X����!q簶s��SO@�Fѩ�e-�DB6D׮z��E$���S�tS�$��뚷!*q�3e�,���_3{�u�JR5a$9���TƁO+x��q\5��
r��Q�K�f]"�,��;A��H�X���/M��5��"���ĩ�/�Z��&�X�'�.㷤��:Tk��dI�>�jü�.��d��<*���R�/�o0���G�I�ru��
߳_F���jl�B�^��cA���.P�J$|����v:'F�n��IC��f|\74�����f�]m�ŭ���U�S��DIF����X����2pŹ=P@��+��+RJ�{����2�*��f�;������G�X��!��q�(� �R�EJ���(Xr߬�C軅f�7>x3��k!֒�Z�iO�\��x`#�τ "�G�'�)$�����5�o!���m�[V\"�9�6�ϐBm��O��&�DdZ4�:@����^p� �8C*�A��b�lj�6ܓa���qq¤�6L�:���C��{E�˿�Մ��c���6*�ݴG���t}&gIʢh�[�&�З�,�����xL�q?�O6:<�\vm-�yp����_^S@�Ui���!�~�%���1&o�9�UL� ���ץz 2��}?�
��2BjB�d�߲��KL[-&M��u�-��R���r<h����j�Gi��X_`>4��h��
�J�2E�Fh�HE%L�"~��F���<(��`H#� �r�������|��t�Q6(�n�������}�/ڨ'���{�P9�ȥ3ӷ��;H��'��\���a)m���h�5�
iE��G�X��Ծ��0�[��[[�Sk2�)ۦfT��Y P�
��)�LX�W������°Pv$��l߸^��|@�)�إ�@�]=�W��p��qE�7PfT� �s"�o��W��곰�����~~S�v���\AD:
��'emc�V�p��ё�r& ��~�ܕUՊ'ggM��g����O���9E|r��go�r��G��B	:���
�؂�nA�p�0�,1�8�{ܖq�Ky����nn�>��'1�2�Or�����c�`�&?���x��0n�G`��U~�UjZ��Z�SN�X�n��<�j�]O6��:��_rS::@D�6�Y��9Fz�i!��G��qI~�cey�Fbt,BDp��m�`�/��(���8E^^���;Χ隩r؉vi�������(Zn�&3���9�l\	���O��!���<��>O?��@�Vdw��:M�J�G_�р����:R��L0Q�}^Z�N����=�p>�l��R��""	���B5�Zr$���[˓��|�.�I��:�R�S��W���rG�'��~�`���Jm�ňz;ͩ��x(:��E��D"ȉk#�u�o�(E�r�p|���Y�u [M�����7�	�v�� <���{}��=�̷x9x��̞����x*m���v����j�`Ы�l�/e���%<�ϠF.���/M:�U��;箤��֛�|j�rr��r7�,��i��m�k��%�FFƹw�4�g-x�B��_�ʔ�2�g��P���UD0�(�r���s��9M����Ӡ�$Q����p�=���y璠�ѱ߅pp�l%M-^(ʎأ�������+�N���VE���(g@���QA?�j����0��$i�u�&����D�,���2YDEm��|��A�'`�����j;��u/���=��ag��뛚� h�P�l�����]��Pa�G�1&��?��M�o��SD�eXF�����e���{i�G=�Ké\X'	�n�{�JL��i*��AP���T֪��+��X�Y�Vc&I��SB:�L�����D2�X�|��>�k�{����Y�o����U��I���;��?����鮅�����_����F�W��]Ok��ٞ(Ӛ��q�'�{ �ю	�;׭�AZ>�<��;�X���X���
^��@�A��ŦY���J|�R����]~ɮ�o]�Nx:��Z�/�`�6Ժc��7��ɇ����.��]���$�:S���t�u0I�a^�f	bϦ�ĆLSǩ�s9n��R+~��Y����L��4X��+�R���i�Yn����i���#|M���#�e\bBo=�������o�`@Or��:�~	�k��GEv�xr�k��[ĝ����@���g�t5 zdE���>�,S�7Fk���x�Ө=�#����V�)b�.h�w�> �!+���!���ը���E��'����{�	�6�R+@g�s┘'�SOTw�ζ ��`\I�գx�H�,���LM2�Ah���H���"�HY�M�^=�U�S�.��T`Į3��߯�B��=?m���6��1�F���VoNkƢ^�=5ͬ��0
_��E�����n�v����E�#�7�/��|����"�Q ��ݜ���6����L�.�q9O�\	�;�=U��2�JU �K�|�y��~=���g.*�Ooҟ��E�R4��6�"�x��9���[Jҗ7CA�q�0+�\"M�6��mKy�x?�Y��g�Z5,Xo߬gCou�vH�#']la���K��ֹ�YEm�B)�Yި�u�N��;����X�5�:T��}�Q(�v�FKCp��똄(�)h9dX��dbB{hYi�B(����'�/����}��Ӻ�L���w���a	i��9s�8:���P��L'��~��/�V��d��ζ�O�ν]�)X�� ���t�d��e�/9��[*$�]��K��a^��m;�3��+F)��-�7 8%$2}B� �����eT�F@K��4.��֐f82�4�(��=�3����5֊ӳB��#���,��^Vr�c��[��n�G����wH�c,}51;r��>51���wx9Q]��(��α�s�5ݭ*�"�ԞK .��	&�������va|��}�o�>;°ϊz�,K����j���A��T��+^]\I-�����7`H|���F�ػ�!6XG?��m��Q�h�s@(��FhM!Ϙ`����=q�-�z��Nr�D�n�c��'b��M�Y��K�kf2�ou:_���.pkԆ�/?p�}����ڴf�xU4�g�
rPy�Ж��no'��+)��*�y}
;��Bd�p��!���:�z��Ǧ�3�c�J�h�H5S����k�c/\N����S����@����@8�0�t�.�l"!'^L��^j��7����{)��u�[�I�,)��~S �9����	Z����$�R�.׉L��+Țpj�����bR����N���MS�A��*ҋP��0�����E�=�.�lX ��n�F����.+�в����� �ϸS��� nX�:�������ۻ�9�J��x� ����_�Ҏ�<ea1([�$T;xH�NW�
���z�R5���nm�#%~|�M�����%�&S�����#�5E�������@�z$H=��0�+FehP�o�E�u��{�O�=ΐ��X�{�t�e�`"��X������ƴ��ݐ��H�F��..�˫�2b�Û��:(M6���Ġ��g��lZ����b�9[�����n��U�g;���H�J��^��(���r�ˇ�ns8 �Q���	S�j����bg���fU�*��Ho��Q�3}��0��fT�hJ�5�En�aØ��=4������"��*<��v.΍��435�������77g�����pm����n���AƱy0D]e�'�����k�_����!ޫ۱�:�&.�**��[�x���J���7F����H��/����4�@�D�ʛ�¡����{t"*0S�&��F��/����Oo}�K�0Y����'b�>]�b���<@�f4=!"��
#�	)Qr�\����&G�5��J�hr |�C�Orp���x�)YZI�Z�,�[M������*1�I��m���w^<�ݨJr�=�s+򘏢�ˋ� D�,����\(%T�g�C%#0m��N����@${#��So����_Q'!G3��&�����_��8pFј56"���<��2���Æ�&dn?PjN	P�FuS�ʭw,�@+gL��}R��P.m���q��6N�~�݁A�>�j	��	�t���ԏy�����*��j�՘_g�	�VsJ����&-(fF;�j�oV��{  �T�<���bu!q)�	U��Q���/q�"�Q����Y�\��̨U��SJ���a����C-bmD^���������:��r<u��fa�P$;�hх�� r��p�س��ٛ�w�����UB���*l�����@�P]���B-���911���{��|?ے���"�{�� �V_�n�+�,7���?S�|G.�c������$ɣ���}HO
㎌w/������<�:n�dц�)���{�ֱY�*�K�+�k�c�b����9?��T93u�����dQsd���M�C�"j>��H@���	~�'���=S×�?�b={�@L�G��:i�,����a�1U�2P�9u�D��Q2x	�C�����C/�	v����OI4?�C9�|�$Pao���w.Lׅl��-�*�vT�
U�E$b�\s�&Y�e�1l�o|��GF����y��'9���۫%
�3��fW�Y�#����i�J�Ҥ�-�:�҂�a.�'�#d������#ї�:v�����AU�@󤸫�c6-�)g{VE��W�SaQ�={�����Mn6 ��uȾH���E�*�~@��r�ź2�x����^%���'5c㝶�l'�"�Q=W(�Z
'k��|��ߎ]�HV�;ʞ�2�U�[9���S+�a�������J,>�_�4?U��1����&�_x��P/+ QԘSq�� 58OH�����:C���Ao�����B����R��Q�֯�y��Ck?{�c���!Q���+N����F�a���蛒8F�,��E��D�D���s�ٰu�L�������T�Qx�O��Z#	��>�jQi��(	]7�_�E�; �҆���̐";��Pq��k�̤.�� ,�I� ���8������h�vvz&�X47Tk�x���g��AVJk���n��՗C�8�� Ԕ��[��bؓ�}[�)�5�Y�NV2��U��>���`�'r��GW��=���~:�3��_V��tCh�M����2@>��stO�Ѱ�C��'"��ԛ�/O��F��I_[�Qɜ�%��;�uS�Y���4�7'����	�=l˭L�ZG�:]P8F`I 2�ت��5M@$�sJ���!Tα��SMTɱ_HZ�F��Hq/r�4xD��q�tw\̎��w�	86k�b6֕��i9�[���W���.�=�[��*F�v�CV,c�� �	��B�n]��ւ�as"�"I\`��=��׀Y���%1���ğc�:�6	�L[I�@RŊ���F��I���������u�?�$�O��$��\�R�@�!�YWL<1DU�q�F�-WE�U1jAj��Ibw�d����rן��%�C����8��	r�S~W�Z����a<Q��㮀|��,T�a�\v���Ȯ?lv���i�!!��=��'�ա�-��psC��^����4d>��8��ɭG�Є�?�����g��Nj�V=3���Oh��R�M`��=�~���y�8���٤?0B�[K7��֌�͍�������HÒ���_I��j�#U9;�v �j�ԋ<��AP$;����q����n�y%���R�~� f��-(ߛ�ٲmHV���2un[�v%A�/�n<��\�	�z�5j�?8��$�Q���v6µ�����h�R�]��ِ�
�����Bh�Nc��	�pٺ?���Ñ����w�O=��l���뤄xᲾb+aj�n�]
�.p�%r���L��/ƐUe~��#�` A�1Kp���G�mȐ�R��B�yu`6�HE(j	���n�|�;���o�$��x8��H���b����tn���Í��r�����꺬F��+9���A_I�	�N�ɩE��b\� ��]|�\�p�V��
?@P7���2����(MRc�/,+�r���/�Kj`�EkP�W�T�%*a9�.����{�ﾮ�|��~=I��m&n��ɞH��X���Y ��3��q��%��P�݅��`0�%<��݋@���5|������ \}�z}����<����F����xksc�'�g� ��^��t�5���������Ӷ;7t�.R�Y���5M���J!�b��$�S@ ܅y�Rݭ��qO2�����W��R�Zq;1}DLX}�]�f���K���qx޾�7]���|��+������՜����Q�=�I��ƃz0��
Dhh�)ݭ��Z�sV^aʪ.�k��Y<	{=Ց�N9������������>S��S�'���Ӣ�4��qDE�\^�j�O�Z�1p�Mک�HR/EC96x 4-+������T\�}�o�aFbH&m���p������޸R�1�ϝ��"���@��w��7u�ބ�HR	8�<7(*��.�el�?Y����f� V����5 � ��sv��i�T��G��Ww��s2Z�b!�]��[cMY*�C3�d���yV�֞��zD�*9�Wd��JS���='X̕6~ng�eE��e!������\Ǽ��H�c6;�YNu�<���1�@l鼤�I:��N��/��nJ�BU�: ��,�=�?��\I� �~]Uq�1'(k�������u�,��ɚ/N Z�m��5h�_e)}H
�|�qhxfn��@�͟47��{�L�}�������z�7kw��V 3��p���F5i�Q�o˽Xߤ�����dАU�m�EM��z�w?/H_��v�����~���M�QKB�w�) ��1$�%py��!C�($ռX�%�W�|k�y!��1��S�͏d9�c��J���f5٣��ep��C��g�Á�ɣ%yi5�=�.@�N]�K
�b;�$�n�=�-}I��3�e�nJ^���sz%:ͰE�m���|4�!I���qU"�feY�Ք�0�%3N�%c���|��j�		�e% ��U~τ�����(o�m�ǞM�r��W)%W��Pe+��/�J�&T`�Ϥw�U[f�F;`xM:����=�<������= ]_��I��r=�����i]�&���t�M���j,M?`��Wm��������=0|\݊��\s�5��Hn:��v��=C �*Y�]p'�L���l~��tk���dA ��`�!�y���f�6����0�ǎS�w�z�R���J.�e�pSx�*(����]���yj�3��zmo�!���5?�r_TW����O-cT�Xs���󬍓��D���Kxo|�^���N�
���6��n7�r��K�{��d)������I'�]�����������˳�K�����9	�S�W�[���Ǘ� )�fc�٬ ? ?]��w�`��.N��pX�A/!_s�����˦Ю_����Łmu��-��{�^B0B-̣���Y!����ΐ� U�D��l*&����I��X]������a��$����M��d��Z�̛��
�«(��E�����V��z��o)� �}��#%�N��ח�#���?����ļ�B�8��|���P6�����0�/<}d8�S����,C�gܮT]_�uSy4�h�����ѹt���~���ͥ��N�?�v% 0gC��ٷ0D��	Y��i�}&DO8(�pÂ9����S��v�K��	����V���'ȿk4�RA|7�DU6$ ����Ҝ!�,���"�BwĜ����|U��0�Q�:��o��" P�R��tw���P��8���o�|�xs�.Ǡ�
F˒�8# �t�����5W�����٤#��W����F�R%��a����ovI���o��h�"���>����0a~vzC"�S"�hyʺ�K��Uu5^�wn�9�!�zj�Y���BǮ�p�o�t�s�@�?H�
ߪ|6$O��DX:D�/�"����ع���~*�k��3�Mx�e�>��&�{�:v�ì(�G3�afY{q�]���a��,�'x�`���8�A��J��-�?�r�����߈��}Q�F�P.�VFM.<��z,[�Jb�%�~vg��q>NQY+���S�3��o��6�8U\Y��7^�g䦜��Tg�\�lJ�������'����X%{im#�[�^� l��C0L�({Е&�e �h��;����Z���C2�	Ѧ^,Md���9d6���U� YF������=k.�YD�MDO Z����D+� qoW~ǘ�n���+���,aЁ�ْz:�ۥ��R��X5c���?.fj<��#��^��N��V5:��l����?�&a*��)c���O����!���L!s�'����^����:<A����+7�)��~1��%���JO���������iO�4<��A��<�Gj��GzU�1-��υ�V��@�J]z��K�(&�O/�A���pZX��\:�ʾ1�� 0�H���c/�6�b}��Q*�)�Y����(`?��
?��7�G��r򱲹�'���$[�M�w/wN�>Ɵ:�/�Y~0����^P�!�����7����(���K���!J�PF'�J��u�ak�5����ߊ���rxl��T�e��������� ��Vn��&A��1���^so�k�5�V�(�e��w�Rh�^C�����\���v�3ۯ�Gt1@B��|J�kj�$�4��Ӝ@�5u�G�8���z��H���w|x��#���)e���EmT~D��vfh=�K[��1�l��9�?S���Y;��
����(��2L?�؋	����A~6>o�D��j>�(��y2{-�~���$ϸp Z�S��QOڔd�X�|5�O���R���Kz�&��w��z�<�+jW��rz��X�a�i��;����Aβ�n$^�W��,{6��{P����yg$�C�9
]ƻ����OΟ�\k�1�Q6,t�`��́tS,�"�J�Tʋ�mg��#7�F�s]0��f:��j�UC�Z��F�d^�ߌtR����z��g�7���p�R�аd��<c��琉���n��#��;���dJ�>��>?%�*�F@N��^c�R򖐁8�z
e�o���o�&{J�n��1�'&g�&l��y��1�<�j�:����e�G~/K�ʬI���
�pma`~Y�M���(ֶ$m���of��4�ۅ��L^��d|:�CfP�
��z���jwm�g���k�7Z?�xi��Q�e�|L��������DA�T'#�ܛ7y	On=�h�1��R�x�P���e��*�ˣAb�q����B*ޢ������3���k��񞑦(/���l�*�[ǇO3����2��9q��%��΀y��,�efr��E3$<��Z,�;�{Y��mi���0f~�`�	-Βf�Jf�`~L�it
e<\�	Pō����X��:�gd�IK7�*��Ꙉg��R�@S9��}��v!�-�浶�G]	0KՌ'�Xv6U�����ڟ�}�8M�8���!hZo/UȰ	�Z���2%{�R��/�P���&�~��T��Sk��`A��kΥ7P@�w���*��&!�W�~�0��YN{!�.p�sy�y�-E0Aw���K= ���P��*��bE����&��seϬ���(��(�X�ԅ�Ĉ��'���x� l1�r�m$KQ���X�8��Tn�j��s%�pl�i���N�Y� �|�E�dЪ񳾥%1�*%�N ��
Ѳ�5y���x?���m.��RM��7Dp�c�Wx��Õnz~in�`����������.�HѶ��j
�S12��v��*���nz��?��>��ϔ�G�I�WP�ѠB�1o\Rr�Ε��HH�V����$3������g� ����{�H�a6�Kx`f;��SVrx��.�!�>��
���$��}{k��h�ݳqZ�)��!�殅d�ׯu�-�0&0|y0L KY�U�1����U�#h �]��r(��z�M�A������VPn��]�=��Ia�B�o�/šZ撾�}�?k��
k&s�2bS,<���(?C�NɈ�'
:�Dw�k1+�0�o	)o9�0�����hv�e�K�,���!A��l��a8��\nKMGU8�(�a&m>T�����^��?��O�փ��_+�x���Z��<���ӡ8���������p�jH߯dC*�$U�.#{	ӟ��誺���R��J~q�/��������� 
���A�p�B���N�ؚ
�h��)[d﷩!(E��o�ؿ������~2�?y�&�y�y�T��?��:�5AK�0���6K�q
!@�hwL�!i�z���6��}�^a��B�3��l�L�5�5Mԇ��^��d�àw�"=� �����C�L�Aʐ��v����ɧ	��r�!�����F���:��H	��7^JČR���L�]�CʠFc`���Z适srSb^��l')l"��_�%I~8v�b��Ǥ~���: � �{���*���m��ƪ�j@3���7L��H�T�K����-�?׳}t�
0T|�@P�^;�-�����c��TLZ4O\��u���F=��s]��L�K)�]����(I�esx&���&���3Ʋm4f�-���k4G�������T�W��|��t�綑y�m	��#�&CГ���S؜,����W�@G�R `�gT���[277va<n���zI�Ihg�]�Ck8�J�
�q���Q 9��ռ�dI���=-L1�+��`r�f
{ڬY��Ԁe�מF���q�r�N�f'ESaJ�� �:�}�!�=[ ���r��n��hRm�`~���S��AO.��*p#1|�ב�S<f�HAg&�ٙK5�b{j�����2�
��a���j�)��!�پƬ��f�OʌPe͈f�z�_���Z>���WY��M0���7�4p�U瞈�}��^[��3����}�)��$�FN�՗��S��`���������}�4�G#�J�?�o�
Ye4�����a0PY�K�]�HU[UX߭b@�v#x������<0WP|\@9T�� pb$���?��W$	H������������8�$M�=D~�$������J=.�>�^}^$(�#��>ᑠ{5��N�ќ�9��AC>$��E;1�@/���>"u�
���\�d5S�+�;�j��$@2�+�$1j���,K��$�N:U˚-��`���}����!�B+�)�ww�[�jk�������st�������=�pC�7/	�q����蛢3�k���[c���E���?E`��<�6�-h�Y"J�!	�i �7�յV���"�_)�neF߻>:���y�-tf\�.t�4�5g�v�<y�����T����;=QOV�$�Nմ^k�E��M��>�C
ִ��E�2��.�Q�}8���ܞeoN�vV/_���b&�<+<|��f��#���xb�zc_bw��� ��4	�t�Y|��p9A�Tyٳ�-��iz�zW#el�h�ಊl��/�J~6���@��Z/8�M�� � �$ �8dn�F�)xu�9'{[�Ψ���M� �1���CE�7�;n�C&+Ƶr����5J�E!@M:��(f��נ��o�f?Bt�7���W��e1J.�o�+�Y��L�I< '[j������o���y����ݙ��_Գ E�U�޷{8j:F=M�W��X�g�O�-�s�R�����7��(�͚�n����V]:M��Q3
��J�6G!�{���)k��e~��QPy'��w.�˥�{o�|��C.��L�׏��l��:����]�gj��2Xd�>����]�I_ C��6�Z��Q�SB"W��GAM���"`oyK���L��ͩT�C1�2���*8�zB�p�ZcO�Z�E�EjG�)i�;��w�kS�$[Am��/q�!摋��D��F���+B����W�u!G|J72�z3��^�F� �0�Q\|��^�
�P����%��7;��,L�䖨9����E?�������<��7�+������k>��8���W<�7@���q`g_�)��M�/����e��5(�ZɶM�[�/]I�U1H��/��Qv2Ut�(K��&��$�2,�$9�����QC��_ݮ��FP�]ʳ�:�DSÃ|�ʣU��h���</��
��:���"��a_p5��Q��D�c<��a�}���l��E�V
�i����^�k�+�g�_��J��@PT�.�ȅ�_u.��$�y�Z_Ϝn��b{��@���7eD����1N"{L)$�p��H}��	1cnO�1wl���v�lb����i��5ԷE��|t��5}�V ���DU�-m�	��㉃��8�q��d�+m��!�e�|�-�w��@O���;�Z�.��jU�EJ�:;	V&	Ը�,a��ݙ%J���U ^����XF˦�:��8}t]���kg���dc�4� >�i��mF|���j����/�D�f���K��86tt3gVE�SN�,��Ȟ�
AqzZP���zo�tK|s�i�;