// fluid_board_soc.v

// Generated using ACDS version 15.1 193

`timescale 1 ps / 1 ps
module fluid_board_soc (
		output wire [15:0] avalon2fpga_slave_0_s2_writedata,                       //                        avalon2fpga_slave_0_s2.writedata
		output wire        avalon2fpga_slave_0_s2_read,                            //                                              .read
		output wire        avalon2fpga_slave_0_s2_write,                           //                                              .write
		output wire [6:0]  avalon2fpga_slave_0_s2_address,                         //                                              .address
		input  wire        avalon2fpga_slave_0_s2_waitrequest,                     //                                              .waitrequest
		input  wire [15:0] avalon2fpga_slave_0_s2_readdata,                        //                                              .readdata
		output wire        avalon_spi_amc7891_1_conduit_end_sclk,                  //              avalon_spi_amc7891_1_conduit_end.sclk
		output wire        avalon_spi_amc7891_1_conduit_end_cs_n,                  //                                              .cs_n
		output wire        avalon_spi_amc7891_1_conduit_end_sdio,                  //                                              .sdio
		input  wire        avalon_spi_amc7891_1_conduit_end_sdo,                   //                                              .sdo
		input  wire        avalon_spi_max31865_0_conduit_end_0_drdy_n,             //           avalon_spi_max31865_0_conduit_end_0.drdy_n
		output wire        avalon_spi_max31865_0_conduit_end_0_sclk,               //                                              .sclk
		output wire        avalon_spi_max31865_0_conduit_end_0_cs_n,               //                                              .cs_n
		output wire        avalon_spi_max31865_0_conduit_end_0_sdi,                //                                              .sdi
		input  wire        avalon_spi_max31865_0_conduit_end_0_sdo,                //                                              .sdo
		input  wire        avalon_spi_max31865_1_conduit_end_0_drdy_n,             //           avalon_spi_max31865_1_conduit_end_0.drdy_n
		output wire        avalon_spi_max31865_1_conduit_end_0_sclk,               //                                              .sclk
		output wire        avalon_spi_max31865_1_conduit_end_0_cs_n,               //                                              .cs_n
		output wire        avalon_spi_max31865_1_conduit_end_0_sdi,                //                                              .sdi
		input  wire        avalon_spi_max31865_1_conduit_end_0_sdo,                //                                              .sdo
		input  wire        avalon_spi_max31865_2_conduit_end_0_drdy_n,             //           avalon_spi_max31865_2_conduit_end_0.drdy_n
		output wire        avalon_spi_max31865_2_conduit_end_0_sclk,               //                                              .sclk
		output wire        avalon_spi_max31865_2_conduit_end_0_cs_n,               //                                              .cs_n
		output wire        avalon_spi_max31865_2_conduit_end_0_sdi,                //                                              .sdi
		input  wire        avalon_spi_max31865_2_conduit_end_0_sdo,                //                                              .sdo
		input  wire        avalon_spi_max31865_3_conduit_end_0_drdy_n,             //           avalon_spi_max31865_3_conduit_end_0.drdy_n
		output wire        avalon_spi_max31865_3_conduit_end_0_sclk,               //                                              .sclk
		output wire        avalon_spi_max31865_3_conduit_end_0_cs_n,               //                                              .cs_n
		output wire        avalon_spi_max31865_3_conduit_end_0_sdi,                //                                              .sdi
		input  wire        avalon_spi_max31865_3_conduit_end_0_sdo,                //                                              .sdo
		input  wire        avalon_spi_max31865_4_conduit_end_0_drdy_n,             //           avalon_spi_max31865_4_conduit_end_0.drdy_n
		output wire        avalon_spi_max31865_4_conduit_end_0_sclk,               //                                              .sclk
		output wire        avalon_spi_max31865_4_conduit_end_0_cs_n,               //                                              .cs_n
		output wire        avalon_spi_max31865_4_conduit_end_0_sdi,                //                                              .sdi
		input  wire        avalon_spi_max31865_4_conduit_end_0_sdo,                //                                              .sdo
		input  wire        avalon_spi_max31865_5_conduit_end_0_drdy_n,             //           avalon_spi_max31865_5_conduit_end_0.drdy_n
		output wire        avalon_spi_max31865_5_conduit_end_0_sclk,               //                                              .sclk
		output wire        avalon_spi_max31865_5_conduit_end_0_cs_n,               //                                              .cs_n
		output wire        avalon_spi_max31865_5_conduit_end_0_sdi,                //                                              .sdi
		input  wire        avalon_spi_max31865_5_conduit_end_0_sdo,                //                                              .sdo
		output wire [3:0]  axi_lw_slave_register_0_conduit_end_0_wr_strb,          //         axi_lw_slave_register_0_conduit_end_0.wr_strb
		output wire        axi_lw_slave_register_0_conduit_end_0_wr_valid,         //                                              .wr_valid
		output wire [15:0] axi_lw_slave_register_0_conduit_end_0_rd_addr,          //                                              .rd_addr
		input  wire [31:0] axi_lw_slave_register_0_conduit_end_0_rd_data,          //                                              .rd_data
		output wire        axi_lw_slave_register_0_conduit_end_0_rd_valid,         //                                              .rd_valid
		input  wire        axi_lw_slave_register_0_conduit_end_0_rd_ready,         //                                              .rd_ready
		output wire [31:0] axi_lw_slave_register_0_conduit_end_0_wr_data,          //                                              .wr_data
		output wire [15:0] axi_lw_slave_register_0_conduit_end_0_wr_addr,          //                                              .wr_addr
		output wire [31:0] flush_pump_pwm_duty_cycle_external_connection_export,   // flush_pump_pwm_duty_cycle_external_connection.export
		output wire [31:0] flush_pump_pwm_freq_external_connection_export,         //       flush_pump_pwm_freq_external_connection.export
		input  wire        hps_0_uart1_cts,                                        //                                   hps_0_uart1.cts
		input  wire        hps_0_uart1_dsr,                                        //                                              .dsr
		input  wire        hps_0_uart1_dcd,                                        //                                              .dcd
		input  wire        hps_0_uart1_ri,                                         //                                              .ri
		output wire        hps_0_uart1_dtr,                                        //                                              .dtr
		output wire        hps_0_uart1_rts,                                        //                                              .rts
		output wire        hps_0_uart1_out1_n,                                     //                                              .out1_n
		output wire        hps_0_uart1_out2_n,                                     //                                              .out2_n
		input  wire        hps_0_uart1_rxd,                                        //                                              .rxd
		output wire        hps_0_uart1_txd,                                        //                                              .txd
		output wire        hps_io_hps_io_emac0_inst_TX_CLK,                        //                                        hps_io.hps_io_emac0_inst_TX_CLK
		output wire        hps_io_hps_io_emac0_inst_TXD0,                          //                                              .hps_io_emac0_inst_TXD0
		output wire        hps_io_hps_io_emac0_inst_TXD1,                          //                                              .hps_io_emac0_inst_TXD1
		output wire        hps_io_hps_io_emac0_inst_TXD2,                          //                                              .hps_io_emac0_inst_TXD2
		output wire        hps_io_hps_io_emac0_inst_TXD3,                          //                                              .hps_io_emac0_inst_TXD3
		input  wire        hps_io_hps_io_emac0_inst_RXD0,                          //                                              .hps_io_emac0_inst_RXD0
		inout  wire        hps_io_hps_io_emac0_inst_MDIO,                          //                                              .hps_io_emac0_inst_MDIO
		output wire        hps_io_hps_io_emac0_inst_MDC,                           //                                              .hps_io_emac0_inst_MDC
		input  wire        hps_io_hps_io_emac0_inst_RX_CTL,                        //                                              .hps_io_emac0_inst_RX_CTL
		output wire        hps_io_hps_io_emac0_inst_TX_CTL,                        //                                              .hps_io_emac0_inst_TX_CTL
		input  wire        hps_io_hps_io_emac0_inst_RX_CLK,                        //                                              .hps_io_emac0_inst_RX_CLK
		input  wire        hps_io_hps_io_emac0_inst_RXD1,                          //                                              .hps_io_emac0_inst_RXD1
		input  wire        hps_io_hps_io_emac0_inst_RXD2,                          //                                              .hps_io_emac0_inst_RXD2
		input  wire        hps_io_hps_io_emac0_inst_RXD3,                          //                                              .hps_io_emac0_inst_RXD3
		inout  wire        hps_io_hps_io_sdio_inst_CMD,                            //                                              .hps_io_sdio_inst_CMD
		inout  wire        hps_io_hps_io_sdio_inst_D0,                             //                                              .hps_io_sdio_inst_D0
		inout  wire        hps_io_hps_io_sdio_inst_D1,                             //                                              .hps_io_sdio_inst_D1
		inout  wire        hps_io_hps_io_sdio_inst_D4,                             //                                              .hps_io_sdio_inst_D4
		inout  wire        hps_io_hps_io_sdio_inst_D5,                             //                                              .hps_io_sdio_inst_D5
		inout  wire        hps_io_hps_io_sdio_inst_D6,                             //                                              .hps_io_sdio_inst_D6
		inout  wire        hps_io_hps_io_sdio_inst_D7,                             //                                              .hps_io_sdio_inst_D7
		output wire        hps_io_hps_io_sdio_inst_CLK,                            //                                              .hps_io_sdio_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_D2,                             //                                              .hps_io_sdio_inst_D2
		inout  wire        hps_io_hps_io_sdio_inst_D3,                             //                                              .hps_io_sdio_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D0,                             //                                              .hps_io_usb1_inst_D0
		inout  wire        hps_io_hps_io_usb1_inst_D1,                             //                                              .hps_io_usb1_inst_D1
		inout  wire        hps_io_hps_io_usb1_inst_D2,                             //                                              .hps_io_usb1_inst_D2
		inout  wire        hps_io_hps_io_usb1_inst_D3,                             //                                              .hps_io_usb1_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D4,                             //                                              .hps_io_usb1_inst_D4
		inout  wire        hps_io_hps_io_usb1_inst_D5,                             //                                              .hps_io_usb1_inst_D5
		inout  wire        hps_io_hps_io_usb1_inst_D6,                             //                                              .hps_io_usb1_inst_D6
		inout  wire        hps_io_hps_io_usb1_inst_D7,                             //                                              .hps_io_usb1_inst_D7
		input  wire        hps_io_hps_io_usb1_inst_CLK,                            //                                              .hps_io_usb1_inst_CLK
		output wire        hps_io_hps_io_usb1_inst_STP,                            //                                              .hps_io_usb1_inst_STP
		input  wire        hps_io_hps_io_usb1_inst_DIR,                            //                                              .hps_io_usb1_inst_DIR
		input  wire        hps_io_hps_io_usb1_inst_NXT,                            //                                              .hps_io_usb1_inst_NXT
		input  wire        hps_io_hps_io_uart0_inst_RX,                            //                                              .hps_io_uart0_inst_RX
		output wire        hps_io_hps_io_uart0_inst_TX,                            //                                              .hps_io_uart0_inst_TX
		inout  wire        hps_io_hps_io_gpio_inst_GPIO37,                         //                                              .hps_io_gpio_inst_GPIO37
		inout  wire        hps_io_hps_io_gpio_inst_GPIO44,                         //                                              .hps_io_gpio_inst_GPIO44
		inout  wire        hps_io_hps_io_gpio_inst_GPIO59,                         //                                              .hps_io_gpio_inst_GPIO59
		inout  wire        i2c_master_d_conduit_end_sda,                           //                      i2c_master_d_conduit_end.sda
		inout  wire        i2c_master_d_conduit_end_scl,                           //                                              .scl
		inout  wire        i2c_master_f_conduit_end_sda,                           //                      i2c_master_f_conduit_end.sda
		inout  wire        i2c_master_f_conduit_end_scl,                           //                                              .scl
		inout  wire        i2c_master_is1_conduit_end_sda,                         //                    i2c_master_is1_conduit_end.sda
		inout  wire        i2c_master_is1_conduit_end_scl,                         //                                              .scl
		inout  wire        i2c_master_is2_conduit_end_sda,                         //                    i2c_master_is2_conduit_end.sda
		inout  wire        i2c_master_is2_conduit_end_scl,                         //                                              .scl
		inout  wire        i2c_master_is3_conduit_end_sda,                         //                    i2c_master_is3_conduit_end.sda
		inout  wire        i2c_master_is3_conduit_end_scl,                         //                                              .scl
		inout  wire        i2c_master_is4_conduit_end_sda,                         //                    i2c_master_is4_conduit_end.sda
		inout  wire        i2c_master_is4_conduit_end_scl,                         //                                              .scl
		inout  wire        i2c_master_p_conduit_end_sda,                           //                      i2c_master_p_conduit_end.sda
		inout  wire        i2c_master_p_conduit_end_scl,                           //                                              .scl
		output wire [14:0] memory_mem_a,                                           //                                        memory.mem_a
		output wire [2:0]  memory_mem_ba,                                          //                                              .mem_ba
		output wire        memory_mem_ck,                                          //                                              .mem_ck
		output wire        memory_mem_ck_n,                                        //                                              .mem_ck_n
		output wire        memory_mem_cke,                                         //                                              .mem_cke
		output wire        memory_mem_cs_n,                                        //                                              .mem_cs_n
		output wire        memory_mem_ras_n,                                       //                                              .mem_ras_n
		output wire        memory_mem_cas_n,                                       //                                              .mem_cas_n
		output wire        memory_mem_we_n,                                        //                                              .mem_we_n
		output wire        memory_mem_reset_n,                                     //                                              .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                                          //                                              .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                                         //                                              .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                                       //                                              .mem_dqs_n
		output wire        memory_mem_odt,                                         //                                              .mem_odt
		output wire [3:0]  memory_mem_dm,                                          //                                              .mem_dm
		input  wire        memory_oct_rzqin,                                       //                                              .oct_rzqin
		input  wire        nios2_qsys_0_cpu_resetrequest_conduit_cpu_resetrequest, //         nios2_qsys_0_cpu_resetrequest_conduit.cpu_resetrequest
		output wire        nios2_qsys_0_cpu_resetrequest_conduit_cpu_resettaken,   //                                              .cpu_resettaken
		input  wire [14:0] pio_input_external_connection_export,                   //                 pio_input_external_connection.export
		output wire [15:0] pio_output_external_connection_export,                  //                pio_output_external_connection.export
		output wire        pio_reset_nios_external_connection_export,              //            pio_reset_nios_external_connection.export
		output wire [31:0] pio_watchdog_cnt_external_connection_export,            //          pio_watchdog_cnt_external_connection.export
		output wire [31:0] pio_watchdog_freq_external_connection_export,           //         pio_watchdog_freq_external_connection.export
		output wire        pll_0_locked_export,                                    //                                  pll_0_locked.export
		input  wire        pll_0_refclk_clk,                                       //                                  pll_0_refclk.clk
		input  wire        pll_0_reset_reset,                                      //                                   pll_0_reset.reset
		output wire        pll_0_sys_clk_clk,                                      //                                 pll_0_sys_clk.clk
		output wire        pll_0_sys_reset_reset_n,                                //                               pll_0_sys_reset.reset_n
		input  wire        qsys_reset_reset_n                                      //                                    qsys_reset.reset_n
	);

	wire  [31:0] nios2_qsys_0_data_master_readdata;                                       // mm_interconnect_0:nios2_qsys_0_data_master_readdata -> nios2_qsys_0:d_readdata
	wire         nios2_qsys_0_data_master_waitrequest;                                    // mm_interconnect_0:nios2_qsys_0_data_master_waitrequest -> nios2_qsys_0:d_waitrequest
	wire         nios2_qsys_0_data_master_debugaccess;                                    // nios2_qsys_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_0_data_master_debugaccess
	wire  [18:0] nios2_qsys_0_data_master_address;                                        // nios2_qsys_0:d_address -> mm_interconnect_0:nios2_qsys_0_data_master_address
	wire   [3:0] nios2_qsys_0_data_master_byteenable;                                     // nios2_qsys_0:d_byteenable -> mm_interconnect_0:nios2_qsys_0_data_master_byteenable
	wire         nios2_qsys_0_data_master_read;                                           // nios2_qsys_0:d_read -> mm_interconnect_0:nios2_qsys_0_data_master_read
	wire         nios2_qsys_0_data_master_write;                                          // nios2_qsys_0:d_write -> mm_interconnect_0:nios2_qsys_0_data_master_write
	wire  [31:0] nios2_qsys_0_data_master_writedata;                                      // nios2_qsys_0:d_writedata -> mm_interconnect_0:nios2_qsys_0_data_master_writedata
	wire   [1:0] hps_0_h2f_axi_master_awburst;                                            // hps_0:h2f_AWBURST -> mm_interconnect_0:hps_0_h2f_axi_master_awburst
	wire   [3:0] hps_0_h2f_axi_master_arlen;                                              // hps_0:h2f_ARLEN -> mm_interconnect_0:hps_0_h2f_axi_master_arlen
	wire   [7:0] hps_0_h2f_axi_master_wstrb;                                              // hps_0:h2f_WSTRB -> mm_interconnect_0:hps_0_h2f_axi_master_wstrb
	wire         hps_0_h2f_axi_master_wready;                                             // mm_interconnect_0:hps_0_h2f_axi_master_wready -> hps_0:h2f_WREADY
	wire  [11:0] hps_0_h2f_axi_master_rid;                                                // mm_interconnect_0:hps_0_h2f_axi_master_rid -> hps_0:h2f_RID
	wire         hps_0_h2f_axi_master_rready;                                             // hps_0:h2f_RREADY -> mm_interconnect_0:hps_0_h2f_axi_master_rready
	wire   [3:0] hps_0_h2f_axi_master_awlen;                                              // hps_0:h2f_AWLEN -> mm_interconnect_0:hps_0_h2f_axi_master_awlen
	wire  [11:0] hps_0_h2f_axi_master_wid;                                                // hps_0:h2f_WID -> mm_interconnect_0:hps_0_h2f_axi_master_wid
	wire   [3:0] hps_0_h2f_axi_master_arcache;                                            // hps_0:h2f_ARCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_arcache
	wire         hps_0_h2f_axi_master_wvalid;                                             // hps_0:h2f_WVALID -> mm_interconnect_0:hps_0_h2f_axi_master_wvalid
	wire  [29:0] hps_0_h2f_axi_master_araddr;                                             // hps_0:h2f_ARADDR -> mm_interconnect_0:hps_0_h2f_axi_master_araddr
	wire   [2:0] hps_0_h2f_axi_master_arprot;                                             // hps_0:h2f_ARPROT -> mm_interconnect_0:hps_0_h2f_axi_master_arprot
	wire   [2:0] hps_0_h2f_axi_master_awprot;                                             // hps_0:h2f_AWPROT -> mm_interconnect_0:hps_0_h2f_axi_master_awprot
	wire  [63:0] hps_0_h2f_axi_master_wdata;                                              // hps_0:h2f_WDATA -> mm_interconnect_0:hps_0_h2f_axi_master_wdata
	wire         hps_0_h2f_axi_master_arvalid;                                            // hps_0:h2f_ARVALID -> mm_interconnect_0:hps_0_h2f_axi_master_arvalid
	wire   [3:0] hps_0_h2f_axi_master_awcache;                                            // hps_0:h2f_AWCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_awcache
	wire  [11:0] hps_0_h2f_axi_master_arid;                                               // hps_0:h2f_ARID -> mm_interconnect_0:hps_0_h2f_axi_master_arid
	wire   [1:0] hps_0_h2f_axi_master_arlock;                                             // hps_0:h2f_ARLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_arlock
	wire   [1:0] hps_0_h2f_axi_master_awlock;                                             // hps_0:h2f_AWLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_awlock
	wire  [29:0] hps_0_h2f_axi_master_awaddr;                                             // hps_0:h2f_AWADDR -> mm_interconnect_0:hps_0_h2f_axi_master_awaddr
	wire   [1:0] hps_0_h2f_axi_master_bresp;                                              // mm_interconnect_0:hps_0_h2f_axi_master_bresp -> hps_0:h2f_BRESP
	wire         hps_0_h2f_axi_master_arready;                                            // mm_interconnect_0:hps_0_h2f_axi_master_arready -> hps_0:h2f_ARREADY
	wire  [63:0] hps_0_h2f_axi_master_rdata;                                              // mm_interconnect_0:hps_0_h2f_axi_master_rdata -> hps_0:h2f_RDATA
	wire         hps_0_h2f_axi_master_awready;                                            // mm_interconnect_0:hps_0_h2f_axi_master_awready -> hps_0:h2f_AWREADY
	wire   [1:0] hps_0_h2f_axi_master_arburst;                                            // hps_0:h2f_ARBURST -> mm_interconnect_0:hps_0_h2f_axi_master_arburst
	wire   [2:0] hps_0_h2f_axi_master_arsize;                                             // hps_0:h2f_ARSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_arsize
	wire         hps_0_h2f_axi_master_bready;                                             // hps_0:h2f_BREADY -> mm_interconnect_0:hps_0_h2f_axi_master_bready
	wire         hps_0_h2f_axi_master_rlast;                                              // mm_interconnect_0:hps_0_h2f_axi_master_rlast -> hps_0:h2f_RLAST
	wire         hps_0_h2f_axi_master_wlast;                                              // hps_0:h2f_WLAST -> mm_interconnect_0:hps_0_h2f_axi_master_wlast
	wire   [1:0] hps_0_h2f_axi_master_rresp;                                              // mm_interconnect_0:hps_0_h2f_axi_master_rresp -> hps_0:h2f_RRESP
	wire  [11:0] hps_0_h2f_axi_master_awid;                                               // hps_0:h2f_AWID -> mm_interconnect_0:hps_0_h2f_axi_master_awid
	wire  [11:0] hps_0_h2f_axi_master_bid;                                                // mm_interconnect_0:hps_0_h2f_axi_master_bid -> hps_0:h2f_BID
	wire         hps_0_h2f_axi_master_bvalid;                                             // mm_interconnect_0:hps_0_h2f_axi_master_bvalid -> hps_0:h2f_BVALID
	wire   [2:0] hps_0_h2f_axi_master_awsize;                                             // hps_0:h2f_AWSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_awsize
	wire         hps_0_h2f_axi_master_awvalid;                                            // hps_0:h2f_AWVALID -> mm_interconnect_0:hps_0_h2f_axi_master_awvalid
	wire         hps_0_h2f_axi_master_rvalid;                                             // mm_interconnect_0:hps_0_h2f_axi_master_rvalid -> hps_0:h2f_RVALID
	wire  [31:0] fpga_only_master_master_readdata;                                        // mm_interconnect_0:fpga_only_master_master_readdata -> fpga_only_master:master_readdata
	wire         fpga_only_master_master_waitrequest;                                     // mm_interconnect_0:fpga_only_master_master_waitrequest -> fpga_only_master:master_waitrequest
	wire  [31:0] fpga_only_master_master_address;                                         // fpga_only_master:master_address -> mm_interconnect_0:fpga_only_master_master_address
	wire         fpga_only_master_master_read;                                            // fpga_only_master:master_read -> mm_interconnect_0:fpga_only_master_master_read
	wire   [3:0] fpga_only_master_master_byteenable;                                      // fpga_only_master:master_byteenable -> mm_interconnect_0:fpga_only_master_master_byteenable
	wire         fpga_only_master_master_readdatavalid;                                   // mm_interconnect_0:fpga_only_master_master_readdatavalid -> fpga_only_master:master_readdatavalid
	wire         fpga_only_master_master_write;                                           // fpga_only_master:master_write -> mm_interconnect_0:fpga_only_master_master_write
	wire  [31:0] fpga_only_master_master_writedata;                                       // fpga_only_master:master_writedata -> mm_interconnect_0:fpga_only_master_master_writedata
	wire  [31:0] nios2_qsys_0_instruction_master_readdata;                                // mm_interconnect_0:nios2_qsys_0_instruction_master_readdata -> nios2_qsys_0:i_readdata
	wire         nios2_qsys_0_instruction_master_waitrequest;                             // mm_interconnect_0:nios2_qsys_0_instruction_master_waitrequest -> nios2_qsys_0:i_waitrequest
	wire  [16:0] nios2_qsys_0_instruction_master_address;                                 // nios2_qsys_0:i_address -> mm_interconnect_0:nios2_qsys_0_instruction_master_address
	wire         nios2_qsys_0_instruction_master_read;                                    // nios2_qsys_0:i_read -> mm_interconnect_0:nios2_qsys_0_instruction_master_read
	wire         nios2_qsys_0_instruction_master_readdatavalid;                           // mm_interconnect_0:nios2_qsys_0_instruction_master_readdatavalid -> nios2_qsys_0:i_readdatavalid
	wire   [1:0] hps_0_h2f_lw_axi_master_awburst;                                         // hps_0:h2f_lw_AWBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awburst
	wire   [3:0] hps_0_h2f_lw_axi_master_arlen;                                           // hps_0:h2f_lw_ARLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlen
	wire   [3:0] hps_0_h2f_lw_axi_master_wstrb;                                           // hps_0:h2f_lw_WSTRB -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wstrb
	wire         hps_0_h2f_lw_axi_master_wready;                                          // mm_interconnect_0:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire  [11:0] hps_0_h2f_lw_axi_master_rid;                                             // mm_interconnect_0:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire         hps_0_h2f_lw_axi_master_rready;                                          // hps_0:h2f_lw_RREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_rready
	wire   [3:0] hps_0_h2f_lw_axi_master_awlen;                                           // hps_0:h2f_lw_AWLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlen
	wire  [11:0] hps_0_h2f_lw_axi_master_wid;                                             // hps_0:h2f_lw_WID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wid
	wire   [3:0] hps_0_h2f_lw_axi_master_arcache;                                         // hps_0:h2f_lw_ARCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arcache
	wire         hps_0_h2f_lw_axi_master_wvalid;                                          // hps_0:h2f_lw_WVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wvalid
	wire  [20:0] hps_0_h2f_lw_axi_master_araddr;                                          // hps_0:h2f_lw_ARADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_araddr
	wire   [2:0] hps_0_h2f_lw_axi_master_arprot;                                          // hps_0:h2f_lw_ARPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arprot
	wire   [2:0] hps_0_h2f_lw_axi_master_awprot;                                          // hps_0:h2f_lw_AWPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awprot
	wire  [31:0] hps_0_h2f_lw_axi_master_wdata;                                           // hps_0:h2f_lw_WDATA -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wdata
	wire         hps_0_h2f_lw_axi_master_arvalid;                                         // hps_0:h2f_lw_ARVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arvalid
	wire   [3:0] hps_0_h2f_lw_axi_master_awcache;                                         // hps_0:h2f_lw_AWCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awcache
	wire  [11:0] hps_0_h2f_lw_axi_master_arid;                                            // hps_0:h2f_lw_ARID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arid
	wire   [1:0] hps_0_h2f_lw_axi_master_arlock;                                          // hps_0:h2f_lw_ARLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlock
	wire   [1:0] hps_0_h2f_lw_axi_master_awlock;                                          // hps_0:h2f_lw_AWLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlock
	wire  [20:0] hps_0_h2f_lw_axi_master_awaddr;                                          // hps_0:h2f_lw_AWADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awaddr
	wire   [1:0] hps_0_h2f_lw_axi_master_bresp;                                           // mm_interconnect_0:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire         hps_0_h2f_lw_axi_master_arready;                                         // mm_interconnect_0:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire  [31:0] hps_0_h2f_lw_axi_master_rdata;                                           // mm_interconnect_0:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire         hps_0_h2f_lw_axi_master_awready;                                         // mm_interconnect_0:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire   [1:0] hps_0_h2f_lw_axi_master_arburst;                                         // hps_0:h2f_lw_ARBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arburst
	wire   [2:0] hps_0_h2f_lw_axi_master_arsize;                                          // hps_0:h2f_lw_ARSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arsize
	wire         hps_0_h2f_lw_axi_master_bready;                                          // hps_0:h2f_lw_BREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_bready
	wire         hps_0_h2f_lw_axi_master_rlast;                                           // mm_interconnect_0:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire         hps_0_h2f_lw_axi_master_wlast;                                           // hps_0:h2f_lw_WLAST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wlast
	wire   [1:0] hps_0_h2f_lw_axi_master_rresp;                                           // mm_interconnect_0:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire  [11:0] hps_0_h2f_lw_axi_master_awid;                                            // hps_0:h2f_lw_AWID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awid
	wire  [11:0] hps_0_h2f_lw_axi_master_bid;                                             // mm_interconnect_0:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire         hps_0_h2f_lw_axi_master_bvalid;                                          // mm_interconnect_0:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire   [2:0] hps_0_h2f_lw_axi_master_awsize;                                          // hps_0:h2f_lw_AWSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awsize
	wire         hps_0_h2f_lw_axi_master_awvalid;                                         // hps_0:h2f_lw_AWVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awvalid
	wire         hps_0_h2f_lw_axi_master_rvalid;                                          // mm_interconnect_0:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire  [15:0] mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_awaddr;  // mm_interconnect_0:axi_lw_slave_register_0_altera_axi4lite_slave_awaddr -> axi_lw_slave_register_0:axs_awaddr
	wire   [1:0] mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_bresp;   // axi_lw_slave_register_0:axs_bresp -> mm_interconnect_0:axi_lw_slave_register_0_altera_axi4lite_slave_bresp
	wire         mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_arready; // axi_lw_slave_register_0:axs_arready -> mm_interconnect_0:axi_lw_slave_register_0_altera_axi4lite_slave_arready
	wire  [31:0] mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_rdata;   // axi_lw_slave_register_0:axs_rdata -> mm_interconnect_0:axi_lw_slave_register_0_altera_axi4lite_slave_rdata
	wire   [3:0] mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_wstrb;   // mm_interconnect_0:axi_lw_slave_register_0_altera_axi4lite_slave_wstrb -> axi_lw_slave_register_0:axs_wstrb
	wire         mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_wready;  // axi_lw_slave_register_0:axs_wready -> mm_interconnect_0:axi_lw_slave_register_0_altera_axi4lite_slave_wready
	wire         mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_awready; // axi_lw_slave_register_0:axs_awready -> mm_interconnect_0:axi_lw_slave_register_0_altera_axi4lite_slave_awready
	wire         mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_rready;  // mm_interconnect_0:axi_lw_slave_register_0_altera_axi4lite_slave_rready -> axi_lw_slave_register_0:axs_rready
	wire         mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_bready;  // mm_interconnect_0:axi_lw_slave_register_0_altera_axi4lite_slave_bready -> axi_lw_slave_register_0:axs_bready
	wire         mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_wvalid;  // mm_interconnect_0:axi_lw_slave_register_0_altera_axi4lite_slave_wvalid -> axi_lw_slave_register_0:axs_wvalid
	wire  [15:0] mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_araddr;  // mm_interconnect_0:axi_lw_slave_register_0_altera_axi4lite_slave_araddr -> axi_lw_slave_register_0:axs_araddr
	wire   [2:0] mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_arprot;  // mm_interconnect_0:axi_lw_slave_register_0_altera_axi4lite_slave_arprot -> axi_lw_slave_register_0:axs_arprot
	wire   [1:0] mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_rresp;   // axi_lw_slave_register_0:axs_rresp -> mm_interconnect_0:axi_lw_slave_register_0_altera_axi4lite_slave_rresp
	wire   [2:0] mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_awprot;  // mm_interconnect_0:axi_lw_slave_register_0_altera_axi4lite_slave_awprot -> axi_lw_slave_register_0:axs_awprot
	wire  [31:0] mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_wdata;   // mm_interconnect_0:axi_lw_slave_register_0_altera_axi4lite_slave_wdata -> axi_lw_slave_register_0:axs_wdata
	wire         mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_arvalid; // mm_interconnect_0:axi_lw_slave_register_0_altera_axi4lite_slave_arvalid -> axi_lw_slave_register_0:axs_arvalid
	wire         mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_bvalid;  // axi_lw_slave_register_0:axs_bvalid -> mm_interconnect_0:axi_lw_slave_register_0_altera_axi4lite_slave_bvalid
	wire         mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_awvalid; // mm_interconnect_0:axi_lw_slave_register_0_altera_axi4lite_slave_awvalid -> axi_lw_slave_register_0:axs_awvalid
	wire         mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_rvalid;  // axi_lw_slave_register_0:axs_rvalid -> mm_interconnect_0:axi_lw_slave_register_0_altera_axi4lite_slave_rvalid
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;                // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;                  // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;               // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;                   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                      // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;                 // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire         mm_interconnect_0_i2c_master_is1_avalon_slave_chipselect;                // mm_interconnect_0:i2c_master_is1_avalon_slave_chipselect -> i2c_master_is1:wb_stb_i
	wire   [7:0] mm_interconnect_0_i2c_master_is1_avalon_slave_readdata;                  // i2c_master_is1:wb_dat_o -> mm_interconnect_0:i2c_master_is1_avalon_slave_readdata
	wire         mm_interconnect_0_i2c_master_is1_avalon_slave_waitrequest;               // i2c_master_is1:wb_ack_o -> mm_interconnect_0:i2c_master_is1_avalon_slave_waitrequest
	wire   [2:0] mm_interconnect_0_i2c_master_is1_avalon_slave_address;                   // mm_interconnect_0:i2c_master_is1_avalon_slave_address -> i2c_master_is1:wb_adr_i
	wire         mm_interconnect_0_i2c_master_is1_avalon_slave_write;                     // mm_interconnect_0:i2c_master_is1_avalon_slave_write -> i2c_master_is1:wb_we_i
	wire   [7:0] mm_interconnect_0_i2c_master_is1_avalon_slave_writedata;                 // mm_interconnect_0:i2c_master_is1_avalon_slave_writedata -> i2c_master_is1:wb_dat_i
	wire         mm_interconnect_0_i2c_master_is2_avalon_slave_chipselect;                // mm_interconnect_0:i2c_master_is2_avalon_slave_chipselect -> i2c_master_is2:wb_stb_i
	wire   [7:0] mm_interconnect_0_i2c_master_is2_avalon_slave_readdata;                  // i2c_master_is2:wb_dat_o -> mm_interconnect_0:i2c_master_is2_avalon_slave_readdata
	wire         mm_interconnect_0_i2c_master_is2_avalon_slave_waitrequest;               // i2c_master_is2:wb_ack_o -> mm_interconnect_0:i2c_master_is2_avalon_slave_waitrequest
	wire   [2:0] mm_interconnect_0_i2c_master_is2_avalon_slave_address;                   // mm_interconnect_0:i2c_master_is2_avalon_slave_address -> i2c_master_is2:wb_adr_i
	wire         mm_interconnect_0_i2c_master_is2_avalon_slave_write;                     // mm_interconnect_0:i2c_master_is2_avalon_slave_write -> i2c_master_is2:wb_we_i
	wire   [7:0] mm_interconnect_0_i2c_master_is2_avalon_slave_writedata;                 // mm_interconnect_0:i2c_master_is2_avalon_slave_writedata -> i2c_master_is2:wb_dat_i
	wire         mm_interconnect_0_i2c_master_is3_avalon_slave_chipselect;                // mm_interconnect_0:i2c_master_is3_avalon_slave_chipselect -> i2c_master_is3:wb_stb_i
	wire   [7:0] mm_interconnect_0_i2c_master_is3_avalon_slave_readdata;                  // i2c_master_is3:wb_dat_o -> mm_interconnect_0:i2c_master_is3_avalon_slave_readdata
	wire         mm_interconnect_0_i2c_master_is3_avalon_slave_waitrequest;               // i2c_master_is3:wb_ack_o -> mm_interconnect_0:i2c_master_is3_avalon_slave_waitrequest
	wire   [2:0] mm_interconnect_0_i2c_master_is3_avalon_slave_address;                   // mm_interconnect_0:i2c_master_is3_avalon_slave_address -> i2c_master_is3:wb_adr_i
	wire         mm_interconnect_0_i2c_master_is3_avalon_slave_write;                     // mm_interconnect_0:i2c_master_is3_avalon_slave_write -> i2c_master_is3:wb_we_i
	wire   [7:0] mm_interconnect_0_i2c_master_is3_avalon_slave_writedata;                 // mm_interconnect_0:i2c_master_is3_avalon_slave_writedata -> i2c_master_is3:wb_dat_i
	wire         mm_interconnect_0_i2c_master_is4_avalon_slave_chipselect;                // mm_interconnect_0:i2c_master_is4_avalon_slave_chipselect -> i2c_master_is4:wb_stb_i
	wire   [7:0] mm_interconnect_0_i2c_master_is4_avalon_slave_readdata;                  // i2c_master_is4:wb_dat_o -> mm_interconnect_0:i2c_master_is4_avalon_slave_readdata
	wire         mm_interconnect_0_i2c_master_is4_avalon_slave_waitrequest;               // i2c_master_is4:wb_ack_o -> mm_interconnect_0:i2c_master_is4_avalon_slave_waitrequest
	wire   [2:0] mm_interconnect_0_i2c_master_is4_avalon_slave_address;                   // mm_interconnect_0:i2c_master_is4_avalon_slave_address -> i2c_master_is4:wb_adr_i
	wire         mm_interconnect_0_i2c_master_is4_avalon_slave_write;                     // mm_interconnect_0:i2c_master_is4_avalon_slave_write -> i2c_master_is4:wb_we_i
	wire   [7:0] mm_interconnect_0_i2c_master_is4_avalon_slave_writedata;                 // mm_interconnect_0:i2c_master_is4_avalon_slave_writedata -> i2c_master_is4:wb_dat_i
	wire         mm_interconnect_0_i2c_master_p_avalon_slave_chipselect;                  // mm_interconnect_0:i2c_master_p_avalon_slave_chipselect -> i2c_master_p:wb_stb_i
	wire   [7:0] mm_interconnect_0_i2c_master_p_avalon_slave_readdata;                    // i2c_master_p:wb_dat_o -> mm_interconnect_0:i2c_master_p_avalon_slave_readdata
	wire         mm_interconnect_0_i2c_master_p_avalon_slave_waitrequest;                 // i2c_master_p:wb_ack_o -> mm_interconnect_0:i2c_master_p_avalon_slave_waitrequest
	wire   [2:0] mm_interconnect_0_i2c_master_p_avalon_slave_address;                     // mm_interconnect_0:i2c_master_p_avalon_slave_address -> i2c_master_p:wb_adr_i
	wire         mm_interconnect_0_i2c_master_p_avalon_slave_write;                       // mm_interconnect_0:i2c_master_p_avalon_slave_write -> i2c_master_p:wb_we_i
	wire   [7:0] mm_interconnect_0_i2c_master_p_avalon_slave_writedata;                   // mm_interconnect_0:i2c_master_p_avalon_slave_writedata -> i2c_master_p:wb_dat_i
	wire         mm_interconnect_0_i2c_master_f_avalon_slave_chipselect;                  // mm_interconnect_0:i2c_master_f_avalon_slave_chipselect -> i2c_master_f:wb_stb_i
	wire   [7:0] mm_interconnect_0_i2c_master_f_avalon_slave_readdata;                    // i2c_master_f:wb_dat_o -> mm_interconnect_0:i2c_master_f_avalon_slave_readdata
	wire         mm_interconnect_0_i2c_master_f_avalon_slave_waitrequest;                 // i2c_master_f:wb_ack_o -> mm_interconnect_0:i2c_master_f_avalon_slave_waitrequest
	wire   [2:0] mm_interconnect_0_i2c_master_f_avalon_slave_address;                     // mm_interconnect_0:i2c_master_f_avalon_slave_address -> i2c_master_f:wb_adr_i
	wire         mm_interconnect_0_i2c_master_f_avalon_slave_write;                       // mm_interconnect_0:i2c_master_f_avalon_slave_write -> i2c_master_f:wb_we_i
	wire   [7:0] mm_interconnect_0_i2c_master_f_avalon_slave_writedata;                   // mm_interconnect_0:i2c_master_f_avalon_slave_writedata -> i2c_master_f:wb_dat_i
	wire         mm_interconnect_0_i2c_master_d_avalon_slave_chipselect;                  // mm_interconnect_0:i2c_master_d_avalon_slave_chipselect -> i2c_master_d:wb_stb_i
	wire   [7:0] mm_interconnect_0_i2c_master_d_avalon_slave_readdata;                    // i2c_master_d:wb_dat_o -> mm_interconnect_0:i2c_master_d_avalon_slave_readdata
	wire         mm_interconnect_0_i2c_master_d_avalon_slave_waitrequest;                 // i2c_master_d:wb_ack_o -> mm_interconnect_0:i2c_master_d_avalon_slave_waitrequest
	wire   [2:0] mm_interconnect_0_i2c_master_d_avalon_slave_address;                     // mm_interconnect_0:i2c_master_d_avalon_slave_address -> i2c_master_d:wb_adr_i
	wire         mm_interconnect_0_i2c_master_d_avalon_slave_write;                       // mm_interconnect_0:i2c_master_d_avalon_slave_write -> i2c_master_d:wb_we_i
	wire   [7:0] mm_interconnect_0_i2c_master_d_avalon_slave_writedata;                   // mm_interconnect_0:i2c_master_d_avalon_slave_writedata -> i2c_master_d:wb_dat_i
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;                          // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;                           // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_debug_mem_slave_readdata;                 // nios2_qsys_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_qsys_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_qsys_0_debug_mem_slave_waitrequest;              // nios2_qsys_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_qsys_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_qsys_0_debug_mem_slave_debugaccess;              // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_debugaccess -> nios2_qsys_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_qsys_0_debug_mem_slave_address;                  // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_address -> nios2_qsys_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_qsys_0_debug_mem_slave_read;                     // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_read -> nios2_qsys_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_qsys_0_debug_mem_slave_byteenable;               // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_byteenable -> nios2_qsys_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_qsys_0_debug_mem_slave_write;                    // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_write -> nios2_qsys_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_debug_mem_slave_writedata;                // mm_interconnect_0:nios2_qsys_0_debug_mem_slave_writedata -> nios2_qsys_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory_nios_cpu_s1_chipselect;                  // mm_interconnect_0:onchip_memory_nios_cpu_s1_chipselect -> onchip_memory_nios_cpu:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory_nios_cpu_s1_readdata;                    // onchip_memory_nios_cpu:readdata -> mm_interconnect_0:onchip_memory_nios_cpu_s1_readdata
	wire  [13:0] mm_interconnect_0_onchip_memory_nios_cpu_s1_address;                     // mm_interconnect_0:onchip_memory_nios_cpu_s1_address -> onchip_memory_nios_cpu:address
	wire   [3:0] mm_interconnect_0_onchip_memory_nios_cpu_s1_byteenable;                  // mm_interconnect_0:onchip_memory_nios_cpu_s1_byteenable -> onchip_memory_nios_cpu:byteenable
	wire         mm_interconnect_0_onchip_memory_nios_cpu_s1_write;                       // mm_interconnect_0:onchip_memory_nios_cpu_s1_write -> onchip_memory_nios_cpu:write
	wire  [31:0] mm_interconnect_0_onchip_memory_nios_cpu_s1_writedata;                   // mm_interconnect_0:onchip_memory_nios_cpu_s1_writedata -> onchip_memory_nios_cpu:writedata
	wire         mm_interconnect_0_onchip_memory_nios_cpu_s1_clken;                       // mm_interconnect_0:onchip_memory_nios_cpu_s1_clken -> onchip_memory_nios_cpu:clken
	wire         mm_interconnect_0_timer_0_s1_chipselect;                                 // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                                   // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                                    // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                                      // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                                  // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_0_timer_1_s1_chipselect;                                 // mm_interconnect_0:timer_1_s1_chipselect -> timer_1:chipselect
	wire  [15:0] mm_interconnect_0_timer_1_s1_readdata;                                   // timer_1:readdata -> mm_interconnect_0:timer_1_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_1_s1_address;                                    // mm_interconnect_0:timer_1_s1_address -> timer_1:address
	wire         mm_interconnect_0_timer_1_s1_write;                                      // mm_interconnect_0:timer_1_s1_write -> timer_1:write_n
	wire  [15:0] mm_interconnect_0_timer_1_s1_writedata;                                  // mm_interconnect_0:timer_1_s1_writedata -> timer_1:writedata
	wire         mm_interconnect_0_pio_input_s1_chipselect;                               // mm_interconnect_0:pio_input_s1_chipselect -> pio_input:chipselect
	wire  [31:0] mm_interconnect_0_pio_input_s1_readdata;                                 // pio_input:readdata -> mm_interconnect_0:pio_input_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_input_s1_address;                                  // mm_interconnect_0:pio_input_s1_address -> pio_input:address
	wire         mm_interconnect_0_pio_input_s1_write;                                    // mm_interconnect_0:pio_input_s1_write -> pio_input:write_n
	wire  [31:0] mm_interconnect_0_pio_input_s1_writedata;                                // mm_interconnect_0:pio_input_s1_writedata -> pio_input:writedata
	wire         mm_interconnect_0_pio_output_s1_chipselect;                              // mm_interconnect_0:pio_output_s1_chipselect -> pio_output:chipselect
	wire  [31:0] mm_interconnect_0_pio_output_s1_readdata;                                // pio_output:readdata -> mm_interconnect_0:pio_output_s1_readdata
	wire   [2:0] mm_interconnect_0_pio_output_s1_address;                                 // mm_interconnect_0:pio_output_s1_address -> pio_output:address
	wire         mm_interconnect_0_pio_output_s1_write;                                   // mm_interconnect_0:pio_output_s1_write -> pio_output:write_n
	wire  [31:0] mm_interconnect_0_pio_output_s1_writedata;                               // mm_interconnect_0:pio_output_s1_writedata -> pio_output:writedata
	wire         mm_interconnect_0_onchip_memory_nios_arm_s1_chipselect;                  // mm_interconnect_0:onchip_memory_nios_arm_s1_chipselect -> onchip_memory_nios_arm:chipselect
	wire  [15:0] mm_interconnect_0_onchip_memory_nios_arm_s1_readdata;                    // onchip_memory_nios_arm:readdata -> mm_interconnect_0:onchip_memory_nios_arm_s1_readdata
	wire  [13:0] mm_interconnect_0_onchip_memory_nios_arm_s1_address;                     // mm_interconnect_0:onchip_memory_nios_arm_s1_address -> onchip_memory_nios_arm:address
	wire   [1:0] mm_interconnect_0_onchip_memory_nios_arm_s1_byteenable;                  // mm_interconnect_0:onchip_memory_nios_arm_s1_byteenable -> onchip_memory_nios_arm:byteenable
	wire         mm_interconnect_0_onchip_memory_nios_arm_s1_write;                       // mm_interconnect_0:onchip_memory_nios_arm_s1_write -> onchip_memory_nios_arm:write
	wire  [15:0] mm_interconnect_0_onchip_memory_nios_arm_s1_writedata;                   // mm_interconnect_0:onchip_memory_nios_arm_s1_writedata -> onchip_memory_nios_arm:writedata
	wire         mm_interconnect_0_onchip_memory_nios_arm_s1_clken;                       // mm_interconnect_0:onchip_memory_nios_arm_s1_clken -> onchip_memory_nios_arm:clken
	wire   [7:0] mm_interconnect_0_avalon_spi_max31865_1_s1_readdata;                     // avalon_spi_max31865_1:avs_s1_readdata -> mm_interconnect_0:avalon_spi_max31865_1_s1_readdata
	wire         mm_interconnect_0_avalon_spi_max31865_1_s1_waitrequest;                  // avalon_spi_max31865_1:avs_s1_waitrequest -> mm_interconnect_0:avalon_spi_max31865_1_s1_waitrequest
	wire   [3:0] mm_interconnect_0_avalon_spi_max31865_1_s1_address;                      // mm_interconnect_0:avalon_spi_max31865_1_s1_address -> avalon_spi_max31865_1:avs_s1_address
	wire         mm_interconnect_0_avalon_spi_max31865_1_s1_read;                         // mm_interconnect_0:avalon_spi_max31865_1_s1_read -> avalon_spi_max31865_1:avs_s1_read
	wire         mm_interconnect_0_avalon_spi_max31865_1_s1_write;                        // mm_interconnect_0:avalon_spi_max31865_1_s1_write -> avalon_spi_max31865_1:avs_s1_write
	wire   [7:0] mm_interconnect_0_avalon_spi_max31865_1_s1_writedata;                    // mm_interconnect_0:avalon_spi_max31865_1_s1_writedata -> avalon_spi_max31865_1:avs_s1_writedata
	wire   [7:0] mm_interconnect_0_avalon_spi_max31865_2_s1_readdata;                     // avalon_spi_max31865_2:avs_s1_readdata -> mm_interconnect_0:avalon_spi_max31865_2_s1_readdata
	wire         mm_interconnect_0_avalon_spi_max31865_2_s1_waitrequest;                  // avalon_spi_max31865_2:avs_s1_waitrequest -> mm_interconnect_0:avalon_spi_max31865_2_s1_waitrequest
	wire   [3:0] mm_interconnect_0_avalon_spi_max31865_2_s1_address;                      // mm_interconnect_0:avalon_spi_max31865_2_s1_address -> avalon_spi_max31865_2:avs_s1_address
	wire         mm_interconnect_0_avalon_spi_max31865_2_s1_read;                         // mm_interconnect_0:avalon_spi_max31865_2_s1_read -> avalon_spi_max31865_2:avs_s1_read
	wire         mm_interconnect_0_avalon_spi_max31865_2_s1_write;                        // mm_interconnect_0:avalon_spi_max31865_2_s1_write -> avalon_spi_max31865_2:avs_s1_write
	wire   [7:0] mm_interconnect_0_avalon_spi_max31865_2_s1_writedata;                    // mm_interconnect_0:avalon_spi_max31865_2_s1_writedata -> avalon_spi_max31865_2:avs_s1_writedata
	wire   [7:0] mm_interconnect_0_avalon_spi_max31865_3_s1_readdata;                     // avalon_spi_max31865_3:avs_s1_readdata -> mm_interconnect_0:avalon_spi_max31865_3_s1_readdata
	wire         mm_interconnect_0_avalon_spi_max31865_3_s1_waitrequest;                  // avalon_spi_max31865_3:avs_s1_waitrequest -> mm_interconnect_0:avalon_spi_max31865_3_s1_waitrequest
	wire   [3:0] mm_interconnect_0_avalon_spi_max31865_3_s1_address;                      // mm_interconnect_0:avalon_spi_max31865_3_s1_address -> avalon_spi_max31865_3:avs_s1_address
	wire         mm_interconnect_0_avalon_spi_max31865_3_s1_read;                         // mm_interconnect_0:avalon_spi_max31865_3_s1_read -> avalon_spi_max31865_3:avs_s1_read
	wire         mm_interconnect_0_avalon_spi_max31865_3_s1_write;                        // mm_interconnect_0:avalon_spi_max31865_3_s1_write -> avalon_spi_max31865_3:avs_s1_write
	wire   [7:0] mm_interconnect_0_avalon_spi_max31865_3_s1_writedata;                    // mm_interconnect_0:avalon_spi_max31865_3_s1_writedata -> avalon_spi_max31865_3:avs_s1_writedata
	wire   [7:0] mm_interconnect_0_avalon_spi_max31865_4_s1_readdata;                     // avalon_spi_max31865_4:avs_s1_readdata -> mm_interconnect_0:avalon_spi_max31865_4_s1_readdata
	wire         mm_interconnect_0_avalon_spi_max31865_4_s1_waitrequest;                  // avalon_spi_max31865_4:avs_s1_waitrequest -> mm_interconnect_0:avalon_spi_max31865_4_s1_waitrequest
	wire   [3:0] mm_interconnect_0_avalon_spi_max31865_4_s1_address;                      // mm_interconnect_0:avalon_spi_max31865_4_s1_address -> avalon_spi_max31865_4:avs_s1_address
	wire         mm_interconnect_0_avalon_spi_max31865_4_s1_read;                         // mm_interconnect_0:avalon_spi_max31865_4_s1_read -> avalon_spi_max31865_4:avs_s1_read
	wire         mm_interconnect_0_avalon_spi_max31865_4_s1_write;                        // mm_interconnect_0:avalon_spi_max31865_4_s1_write -> avalon_spi_max31865_4:avs_s1_write
	wire   [7:0] mm_interconnect_0_avalon_spi_max31865_4_s1_writedata;                    // mm_interconnect_0:avalon_spi_max31865_4_s1_writedata -> avalon_spi_max31865_4:avs_s1_writedata
	wire   [7:0] mm_interconnect_0_avalon_spi_max31865_5_s1_readdata;                     // avalon_spi_max31865_5:avs_s1_readdata -> mm_interconnect_0:avalon_spi_max31865_5_s1_readdata
	wire         mm_interconnect_0_avalon_spi_max31865_5_s1_waitrequest;                  // avalon_spi_max31865_5:avs_s1_waitrequest -> mm_interconnect_0:avalon_spi_max31865_5_s1_waitrequest
	wire   [3:0] mm_interconnect_0_avalon_spi_max31865_5_s1_address;                      // mm_interconnect_0:avalon_spi_max31865_5_s1_address -> avalon_spi_max31865_5:avs_s1_address
	wire         mm_interconnect_0_avalon_spi_max31865_5_s1_read;                         // mm_interconnect_0:avalon_spi_max31865_5_s1_read -> avalon_spi_max31865_5:avs_s1_read
	wire         mm_interconnect_0_avalon_spi_max31865_5_s1_write;                        // mm_interconnect_0:avalon_spi_max31865_5_s1_write -> avalon_spi_max31865_5:avs_s1_write
	wire   [7:0] mm_interconnect_0_avalon_spi_max31865_5_s1_writedata;                    // mm_interconnect_0:avalon_spi_max31865_5_s1_writedata -> avalon_spi_max31865_5:avs_s1_writedata
	wire   [7:0] mm_interconnect_0_avalon_spi_max31865_0_s1_readdata;                     // avalon_spi_max31865_0:avs_s1_readdata -> mm_interconnect_0:avalon_spi_max31865_0_s1_readdata
	wire         mm_interconnect_0_avalon_spi_max31865_0_s1_waitrequest;                  // avalon_spi_max31865_0:avs_s1_waitrequest -> mm_interconnect_0:avalon_spi_max31865_0_s1_waitrequest
	wire   [3:0] mm_interconnect_0_avalon_spi_max31865_0_s1_address;                      // mm_interconnect_0:avalon_spi_max31865_0_s1_address -> avalon_spi_max31865_0:avs_s1_address
	wire         mm_interconnect_0_avalon_spi_max31865_0_s1_read;                         // mm_interconnect_0:avalon_spi_max31865_0_s1_read -> avalon_spi_max31865_0:avs_s1_read
	wire         mm_interconnect_0_avalon_spi_max31865_0_s1_write;                        // mm_interconnect_0:avalon_spi_max31865_0_s1_write -> avalon_spi_max31865_0:avs_s1_write
	wire   [7:0] mm_interconnect_0_avalon_spi_max31865_0_s1_writedata;                    // mm_interconnect_0:avalon_spi_max31865_0_s1_writedata -> avalon_spi_max31865_0:avs_s1_writedata
	wire  [15:0] mm_interconnect_0_avalon_spi_amc7891_1_s1_readdata;                      // avalon_spi_amc7891_1:avs_s1_readdata -> mm_interconnect_0:avalon_spi_amc7891_1_s1_readdata
	wire         mm_interconnect_0_avalon_spi_amc7891_1_s1_waitrequest;                   // avalon_spi_amc7891_1:avs_s1_waitrequest -> mm_interconnect_0:avalon_spi_amc7891_1_s1_waitrequest
	wire   [6:0] mm_interconnect_0_avalon_spi_amc7891_1_s1_address;                       // mm_interconnect_0:avalon_spi_amc7891_1_s1_address -> avalon_spi_amc7891_1:avs_s1_address
	wire         mm_interconnect_0_avalon_spi_amc7891_1_s1_read;                          // mm_interconnect_0:avalon_spi_amc7891_1_s1_read -> avalon_spi_amc7891_1:avs_s1_read
	wire         mm_interconnect_0_avalon_spi_amc7891_1_s1_write;                         // mm_interconnect_0:avalon_spi_amc7891_1_s1_write -> avalon_spi_amc7891_1:avs_s1_write
	wire  [15:0] mm_interconnect_0_avalon_spi_amc7891_1_s1_writedata;                     // mm_interconnect_0:avalon_spi_amc7891_1_s1_writedata -> avalon_spi_amc7891_1:avs_s1_writedata
	wire         mm_interconnect_0_flush_pump_pwm_duty_cycle_s1_chipselect;               // mm_interconnect_0:flush_pump_pwm_duty_cycle_s1_chipselect -> flush_pump_pwm_duty_cycle:chipselect
	wire  [31:0] mm_interconnect_0_flush_pump_pwm_duty_cycle_s1_readdata;                 // flush_pump_pwm_duty_cycle:readdata -> mm_interconnect_0:flush_pump_pwm_duty_cycle_s1_readdata
	wire   [1:0] mm_interconnect_0_flush_pump_pwm_duty_cycle_s1_address;                  // mm_interconnect_0:flush_pump_pwm_duty_cycle_s1_address -> flush_pump_pwm_duty_cycle:address
	wire         mm_interconnect_0_flush_pump_pwm_duty_cycle_s1_write;                    // mm_interconnect_0:flush_pump_pwm_duty_cycle_s1_write -> flush_pump_pwm_duty_cycle:write_n
	wire  [31:0] mm_interconnect_0_flush_pump_pwm_duty_cycle_s1_writedata;                // mm_interconnect_0:flush_pump_pwm_duty_cycle_s1_writedata -> flush_pump_pwm_duty_cycle:writedata
	wire         mm_interconnect_0_flush_pump_pwm_freq_s1_chipselect;                     // mm_interconnect_0:flush_pump_pwm_freq_s1_chipselect -> flush_pump_pwm_freq:chipselect
	wire  [31:0] mm_interconnect_0_flush_pump_pwm_freq_s1_readdata;                       // flush_pump_pwm_freq:readdata -> mm_interconnect_0:flush_pump_pwm_freq_s1_readdata
	wire   [1:0] mm_interconnect_0_flush_pump_pwm_freq_s1_address;                        // mm_interconnect_0:flush_pump_pwm_freq_s1_address -> flush_pump_pwm_freq:address
	wire         mm_interconnect_0_flush_pump_pwm_freq_s1_write;                          // mm_interconnect_0:flush_pump_pwm_freq_s1_write -> flush_pump_pwm_freq:write_n
	wire  [31:0] mm_interconnect_0_flush_pump_pwm_freq_s1_writedata;                      // mm_interconnect_0:flush_pump_pwm_freq_s1_writedata -> flush_pump_pwm_freq:writedata
	wire         mm_interconnect_0_timer_2_s1_chipselect;                                 // mm_interconnect_0:timer_2_s1_chipselect -> timer_2:chipselect
	wire  [15:0] mm_interconnect_0_timer_2_s1_readdata;                                   // timer_2:readdata -> mm_interconnect_0:timer_2_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_2_s1_address;                                    // mm_interconnect_0:timer_2_s1_address -> timer_2:address
	wire         mm_interconnect_0_timer_2_s1_write;                                      // mm_interconnect_0:timer_2_s1_write -> timer_2:write_n
	wire  [15:0] mm_interconnect_0_timer_2_s1_writedata;                                  // mm_interconnect_0:timer_2_s1_writedata -> timer_2:writedata
	wire         mm_interconnect_0_pio_watchdog_freq_s1_chipselect;                       // mm_interconnect_0:pio_watchdog_freq_s1_chipselect -> pio_watchdog_freq:chipselect
	wire  [31:0] mm_interconnect_0_pio_watchdog_freq_s1_readdata;                         // pio_watchdog_freq:readdata -> mm_interconnect_0:pio_watchdog_freq_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_watchdog_freq_s1_address;                          // mm_interconnect_0:pio_watchdog_freq_s1_address -> pio_watchdog_freq:address
	wire         mm_interconnect_0_pio_watchdog_freq_s1_write;                            // mm_interconnect_0:pio_watchdog_freq_s1_write -> pio_watchdog_freq:write_n
	wire  [31:0] mm_interconnect_0_pio_watchdog_freq_s1_writedata;                        // mm_interconnect_0:pio_watchdog_freq_s1_writedata -> pio_watchdog_freq:writedata
	wire         mm_interconnect_0_pio_watchdog_cnt_s1_chipselect;                        // mm_interconnect_0:pio_watchdog_cnt_s1_chipselect -> pio_watchdog_cnt:chipselect
	wire  [31:0] mm_interconnect_0_pio_watchdog_cnt_s1_readdata;                          // pio_watchdog_cnt:readdata -> mm_interconnect_0:pio_watchdog_cnt_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_watchdog_cnt_s1_address;                           // mm_interconnect_0:pio_watchdog_cnt_s1_address -> pio_watchdog_cnt:address
	wire         mm_interconnect_0_pio_watchdog_cnt_s1_write;                             // mm_interconnect_0:pio_watchdog_cnt_s1_write -> pio_watchdog_cnt:write_n
	wire  [31:0] mm_interconnect_0_pio_watchdog_cnt_s1_writedata;                         // mm_interconnect_0:pio_watchdog_cnt_s1_writedata -> pio_watchdog_cnt:writedata
	wire  [15:0] mm_interconnect_0_avalon2fpga_slave_0_s1_readdata;                       // avalon2fpga_slave_0:avs_s1_readdata -> mm_interconnect_0:avalon2fpga_slave_0_s1_readdata
	wire         mm_interconnect_0_avalon2fpga_slave_0_s1_waitrequest;                    // avalon2fpga_slave_0:avs_s1_waitrequest -> mm_interconnect_0:avalon2fpga_slave_0_s1_waitrequest
	wire   [6:0] mm_interconnect_0_avalon2fpga_slave_0_s1_address;                        // mm_interconnect_0:avalon2fpga_slave_0_s1_address -> avalon2fpga_slave_0:avs_s1_address
	wire         mm_interconnect_0_avalon2fpga_slave_0_s1_read;                           // mm_interconnect_0:avalon2fpga_slave_0_s1_read -> avalon2fpga_slave_0:avs_s1_read
	wire         mm_interconnect_0_avalon2fpga_slave_0_s1_write;                          // mm_interconnect_0:avalon2fpga_slave_0_s1_write -> avalon2fpga_slave_0:avs_s1_write
	wire  [15:0] mm_interconnect_0_avalon2fpga_slave_0_s1_writedata;                      // mm_interconnect_0:avalon2fpga_slave_0_s1_writedata -> avalon2fpga_slave_0:avs_s1_writedata
	wire         mm_interconnect_0_onchip_memory_nios_cpu_s2_chipselect;                  // mm_interconnect_0:onchip_memory_nios_cpu_s2_chipselect -> onchip_memory_nios_cpu:chipselect2
	wire  [31:0] mm_interconnect_0_onchip_memory_nios_cpu_s2_readdata;                    // onchip_memory_nios_cpu:readdata2 -> mm_interconnect_0:onchip_memory_nios_cpu_s2_readdata
	wire  [13:0] mm_interconnect_0_onchip_memory_nios_cpu_s2_address;                     // mm_interconnect_0:onchip_memory_nios_cpu_s2_address -> onchip_memory_nios_cpu:address2
	wire   [3:0] mm_interconnect_0_onchip_memory_nios_cpu_s2_byteenable;                  // mm_interconnect_0:onchip_memory_nios_cpu_s2_byteenable -> onchip_memory_nios_cpu:byteenable2
	wire         mm_interconnect_0_onchip_memory_nios_cpu_s2_write;                       // mm_interconnect_0:onchip_memory_nios_cpu_s2_write -> onchip_memory_nios_cpu:write2
	wire  [31:0] mm_interconnect_0_onchip_memory_nios_cpu_s2_writedata;                   // mm_interconnect_0:onchip_memory_nios_cpu_s2_writedata -> onchip_memory_nios_cpu:writedata2
	wire         mm_interconnect_0_onchip_memory_nios_cpu_s2_clken;                       // mm_interconnect_0:onchip_memory_nios_cpu_s2_clken -> onchip_memory_nios_cpu:clken2
	wire         mm_interconnect_0_onchip_memory_nios_arm_s2_chipselect;                  // mm_interconnect_0:onchip_memory_nios_arm_s2_chipselect -> onchip_memory_nios_arm:chipselect2
	wire  [15:0] mm_interconnect_0_onchip_memory_nios_arm_s2_readdata;                    // onchip_memory_nios_arm:readdata2 -> mm_interconnect_0:onchip_memory_nios_arm_s2_readdata
	wire  [13:0] mm_interconnect_0_onchip_memory_nios_arm_s2_address;                     // mm_interconnect_0:onchip_memory_nios_arm_s2_address -> onchip_memory_nios_arm:address2
	wire   [1:0] mm_interconnect_0_onchip_memory_nios_arm_s2_byteenable;                  // mm_interconnect_0:onchip_memory_nios_arm_s2_byteenable -> onchip_memory_nios_arm:byteenable2
	wire         mm_interconnect_0_onchip_memory_nios_arm_s2_write;                       // mm_interconnect_0:onchip_memory_nios_arm_s2_write -> onchip_memory_nios_arm:write2
	wire  [15:0] mm_interconnect_0_onchip_memory_nios_arm_s2_writedata;                   // mm_interconnect_0:onchip_memory_nios_arm_s2_writedata -> onchip_memory_nios_arm:writedata2
	wire         mm_interconnect_0_onchip_memory_nios_arm_s2_clken;                       // mm_interconnect_0:onchip_memory_nios_arm_s2_clken -> onchip_memory_nios_arm:clken2
	wire         mm_interconnect_0_pio_reset_nios_s1_chipselect;                          // mm_interconnect_0:pio_reset_nios_s1_chipselect -> pio_reset_nios:chipselect
	wire  [31:0] mm_interconnect_0_pio_reset_nios_s1_readdata;                            // pio_reset_nios:readdata -> mm_interconnect_0:pio_reset_nios_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_reset_nios_s1_address;                             // mm_interconnect_0:pio_reset_nios_s1_address -> pio_reset_nios:address
	wire         mm_interconnect_0_pio_reset_nios_s1_write;                               // mm_interconnect_0:pio_reset_nios_s1_write -> pio_reset_nios:write_n
	wire  [31:0] mm_interconnect_0_pio_reset_nios_s1_writedata;                           // mm_interconnect_0:pio_reset_nios_s1_writedata -> pio_reset_nios:writedata
	wire  [31:0] hps_0_f2h_irq0_irq;                                                      // irq_mapper:sender_irq -> hps_0:f2h_irq_p0
	wire  [31:0] hps_0_f2h_irq1_irq;                                                      // irq_mapper_001:sender_irq -> hps_0:f2h_irq_p1
	wire         irq_mapper_002_receiver0_irq;                                            // i2c_master_is1:wb_inta_o -> irq_mapper_002:receiver0_irq
	wire         irq_mapper_002_receiver1_irq;                                            // i2c_master_is2:wb_inta_o -> irq_mapper_002:receiver1_irq
	wire         irq_mapper_002_receiver2_irq;                                            // i2c_master_is3:wb_inta_o -> irq_mapper_002:receiver2_irq
	wire         irq_mapper_002_receiver3_irq;                                            // i2c_master_is4:wb_inta_o -> irq_mapper_002:receiver3_irq
	wire         irq_mapper_002_receiver4_irq;                                            // i2c_master_p:wb_inta_o -> irq_mapper_002:receiver4_irq
	wire         irq_mapper_002_receiver5_irq;                                            // i2c_master_f:wb_inta_o -> irq_mapper_002:receiver5_irq
	wire         irq_mapper_002_receiver6_irq;                                            // i2c_master_d:wb_inta_o -> irq_mapper_002:receiver6_irq
	wire         irq_mapper_002_receiver7_irq;                                            // timer_0:irq -> irq_mapper_002:receiver7_irq
	wire         irq_mapper_002_receiver8_irq;                                            // timer_1:irq -> irq_mapper_002:receiver8_irq
	wire         irq_mapper_002_receiver9_irq;                                            // pio_input:irq -> irq_mapper_002:receiver9_irq
	wire         irq_mapper_002_receiver11_irq;                                           // timer_2:irq -> irq_mapper_002:receiver11_irq
	wire  [31:0] nios2_qsys_0_irq_irq;                                                    // irq_mapper_002:sender_irq -> nios2_qsys_0:irq
	wire         irq_mapper_receiver0_irq;                                                // jtag_uart:av_irq -> [irq_mapper:receiver0_irq, irq_mapper_002:receiver10_irq]
	wire         rst_controller_reset_out_reset;                                          // rst_controller:reset_out -> [avalon2fpga_slave_0:rsi_reset_reset_n, avalon_spi_amc7891_1:csi_clock_reset_n, avalon_spi_max31865_0:rsi_reset_reset_n, avalon_spi_max31865_1:rsi_reset_reset_n, avalon_spi_max31865_2:rsi_reset_reset_n, avalon_spi_max31865_3:rsi_reset_reset_n, avalon_spi_max31865_4:rsi_reset_reset_n, avalon_spi_max31865_5:rsi_reset_reset_n, axi_lw_slave_register_0:rsi_reset_reset_n, flush_pump_pwm_duty_cycle:reset_n, flush_pump_pwm_freq:reset_n, i2c_master_d:wb_rst_i, i2c_master_f:wb_rst_i, i2c_master_is1:wb_rst_i, i2c_master_is2:wb_rst_i, i2c_master_is3:wb_rst_i, i2c_master_is4:wb_rst_i, i2c_master_p:wb_rst_i, irq_mapper_002:reset, jtag_uart:rst_n, mm_interconnect_0:fpga_only_master_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_0:nios2_qsys_0_reset_reset_bridge_in_reset_reset, nios2_qsys_0:reset_n, pio_input:reset_n, pio_output:reset_n, pio_watchdog_cnt:reset_n, pio_watchdog_freq:reset_n, rst_translator:in_reset, timer_0:reset_n, timer_1:reset_n, timer_2:reset_n]
	wire         rst_controller_reset_out_reset_req;                                      // rst_controller:reset_req -> [nios2_qsys_0:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                                      // rst_controller_001:reset_out -> [mm_interconnect_0:sysid_reset_reset_bridge_in_reset_reset, onchip_memory_nios_arm:reset, onchip_memory_nios_cpu:reset, pio_reset_nios:reset_n, rst_translator_001:in_reset, sysid:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                                  // rst_controller_001:reset_req -> [onchip_memory_nios_arm:reset_req, onchip_memory_nios_cpu:reset_req, rst_translator_001:reset_req_in]
	wire         hps_0_h2f_reset_reset;                                                   // hps_0:h2f_rst_n -> [rst_controller_001:reset_in1, rst_controller_002:reset_in0]
	wire         rst_controller_002_reset_out_reset;                                      // rst_controller_002:reset_out -> mm_interconnect_0:hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset

	avalon2fpga_slave #(
		.g_address_width (7),
		.g_data_width    (16)
	) avalon2fpga_slave_0 (
		.csi_clock_clk      (pll_0_sys_clk_clk),                                    // clock.clk
		.rsi_reset_reset_n  (~rst_controller_reset_out_reset),                      // reset.reset_n
		.avs_s1_writedata   (mm_interconnect_0_avalon2fpga_slave_0_s1_writedata),   //    s1.writedata
		.avs_s1_read        (mm_interconnect_0_avalon2fpga_slave_0_s1_read),        //      .read
		.avs_s1_write       (mm_interconnect_0_avalon2fpga_slave_0_s1_write),       //      .write
		.avs_s1_address     (mm_interconnect_0_avalon2fpga_slave_0_s1_address),     //      .address
		.avs_s1_waitrequest (mm_interconnect_0_avalon2fpga_slave_0_s1_waitrequest), //      .waitrequest
		.avs_s1_readdata    (mm_interconnect_0_avalon2fpga_slave_0_s1_readdata),    //      .readdata
		.avm_s2_writedata   (avalon2fpga_slave_0_s2_writedata),                     //    s2.writedata
		.avm_s2_read        (avalon2fpga_slave_0_s2_read),                          //      .read
		.avm_s2_write       (avalon2fpga_slave_0_s2_write),                         //      .write
		.avm_s2_address     (avalon2fpga_slave_0_s2_address),                       //      .address
		.avm_s2_waitrequest (avalon2fpga_slave_0_s2_waitrequest),                   //      .waitrequest
		.avm_s2_readdata    (avalon2fpga_slave_0_s2_readdata)                       //      .readdata
	);

	avalon_spi_AMC7891 avalon_spi_amc7891_1 (
		.csi_clock_clk      (pll_0_sys_clk_clk),                                     //       clock.clk
		.csi_clock_reset_n  (~rst_controller_reset_out_reset),                       // clock_reset.reset_n
		.avs_s1_writedata   (mm_interconnect_0_avalon_spi_amc7891_1_s1_writedata),   //          s1.writedata
		.avs_s1_read        (mm_interconnect_0_avalon_spi_amc7891_1_s1_read),        //            .read
		.avs_s1_write       (mm_interconnect_0_avalon_spi_amc7891_1_s1_write),       //            .write
		.avs_s1_address     (mm_interconnect_0_avalon_spi_amc7891_1_s1_address),     //            .address
		.avs_s1_waitrequest (mm_interconnect_0_avalon_spi_amc7891_1_s1_waitrequest), //            .waitrequest
		.avs_s1_readdata    (mm_interconnect_0_avalon_spi_amc7891_1_s1_readdata),    //            .readdata
		.coe_s1_sclk        (avalon_spi_amc7891_1_conduit_end_sclk),                 // conduit_end.sclk
		.coe_s1_cs_n        (avalon_spi_amc7891_1_conduit_end_cs_n),                 //            .cs_n
		.coe_s1_sdio        (avalon_spi_amc7891_1_conduit_end_sdio),                 //            .sdio
		.coe_s1_sdo         (avalon_spi_amc7891_1_conduit_end_sdo)                   //            .sdo
	);

	avalon_spi_max31865 #(
		.g_cpol ("'0'")
	) avalon_spi_max31865_0 (
		.csi_clock_clk      (pll_0_sys_clk_clk),                                      //         clock.clk
		.rsi_reset_reset_n  (~rst_controller_reset_out_reset),                        //         reset.reset_n
		.avs_s1_writedata   (mm_interconnect_0_avalon_spi_max31865_0_s1_writedata),   //            s1.writedata
		.avs_s1_read        (mm_interconnect_0_avalon_spi_max31865_0_s1_read),        //              .read
		.avs_s1_write       (mm_interconnect_0_avalon_spi_max31865_0_s1_write),       //              .write
		.avs_s1_address     (mm_interconnect_0_avalon_spi_max31865_0_s1_address),     //              .address
		.avs_s1_waitrequest (mm_interconnect_0_avalon_spi_max31865_0_s1_waitrequest), //              .waitrequest
		.avs_s1_readdata    (mm_interconnect_0_avalon_spi_max31865_0_s1_readdata),    //              .readdata
		.coe_s2_drdy_n      (avalon_spi_max31865_0_conduit_end_0_drdy_n),             // conduit_end_0.drdy_n
		.coe_s2_sclk        (avalon_spi_max31865_0_conduit_end_0_sclk),               //              .sclk
		.coe_s2_cs_n        (avalon_spi_max31865_0_conduit_end_0_cs_n),               //              .cs_n
		.coe_s2_sdi         (avalon_spi_max31865_0_conduit_end_0_sdi),                //              .sdi
		.coe_s2_sdo         (avalon_spi_max31865_0_conduit_end_0_sdo)                 //              .sdo
	);

	avalon_spi_max31865 #(
		.g_cpol ("'0'")
	) avalon_spi_max31865_1 (
		.csi_clock_clk      (pll_0_sys_clk_clk),                                      //         clock.clk
		.rsi_reset_reset_n  (~rst_controller_reset_out_reset),                        //         reset.reset_n
		.avs_s1_writedata   (mm_interconnect_0_avalon_spi_max31865_1_s1_writedata),   //            s1.writedata
		.avs_s1_read        (mm_interconnect_0_avalon_spi_max31865_1_s1_read),        //              .read
		.avs_s1_write       (mm_interconnect_0_avalon_spi_max31865_1_s1_write),       //              .write
		.avs_s1_address     (mm_interconnect_0_avalon_spi_max31865_1_s1_address),     //              .address
		.avs_s1_waitrequest (mm_interconnect_0_avalon_spi_max31865_1_s1_waitrequest), //              .waitrequest
		.avs_s1_readdata    (mm_interconnect_0_avalon_spi_max31865_1_s1_readdata),    //              .readdata
		.coe_s2_drdy_n      (avalon_spi_max31865_1_conduit_end_0_drdy_n),             // conduit_end_0.drdy_n
		.coe_s2_sclk        (avalon_spi_max31865_1_conduit_end_0_sclk),               //              .sclk
		.coe_s2_cs_n        (avalon_spi_max31865_1_conduit_end_0_cs_n),               //              .cs_n
		.coe_s2_sdi         (avalon_spi_max31865_1_conduit_end_0_sdi),                //              .sdi
		.coe_s2_sdo         (avalon_spi_max31865_1_conduit_end_0_sdo)                 //              .sdo
	);

	avalon_spi_max31865 #(
		.g_cpol ("'0'")
	) avalon_spi_max31865_2 (
		.csi_clock_clk      (pll_0_sys_clk_clk),                                      //         clock.clk
		.rsi_reset_reset_n  (~rst_controller_reset_out_reset),                        //         reset.reset_n
		.avs_s1_writedata   (mm_interconnect_0_avalon_spi_max31865_2_s1_writedata),   //            s1.writedata
		.avs_s1_read        (mm_interconnect_0_avalon_spi_max31865_2_s1_read),        //              .read
		.avs_s1_write       (mm_interconnect_0_avalon_spi_max31865_2_s1_write),       //              .write
		.avs_s1_address     (mm_interconnect_0_avalon_spi_max31865_2_s1_address),     //              .address
		.avs_s1_waitrequest (mm_interconnect_0_avalon_spi_max31865_2_s1_waitrequest), //              .waitrequest
		.avs_s1_readdata    (mm_interconnect_0_avalon_spi_max31865_2_s1_readdata),    //              .readdata
		.coe_s2_drdy_n      (avalon_spi_max31865_2_conduit_end_0_drdy_n),             // conduit_end_0.drdy_n
		.coe_s2_sclk        (avalon_spi_max31865_2_conduit_end_0_sclk),               //              .sclk
		.coe_s2_cs_n        (avalon_spi_max31865_2_conduit_end_0_cs_n),               //              .cs_n
		.coe_s2_sdi         (avalon_spi_max31865_2_conduit_end_0_sdi),                //              .sdi
		.coe_s2_sdo         (avalon_spi_max31865_2_conduit_end_0_sdo)                 //              .sdo
	);

	avalon_spi_max31865 #(
		.g_cpol ("'0'")
	) avalon_spi_max31865_3 (
		.csi_clock_clk      (pll_0_sys_clk_clk),                                      //         clock.clk
		.rsi_reset_reset_n  (~rst_controller_reset_out_reset),                        //         reset.reset_n
		.avs_s1_writedata   (mm_interconnect_0_avalon_spi_max31865_3_s1_writedata),   //            s1.writedata
		.avs_s1_read        (mm_interconnect_0_avalon_spi_max31865_3_s1_read),        //              .read
		.avs_s1_write       (mm_interconnect_0_avalon_spi_max31865_3_s1_write),       //              .write
		.avs_s1_address     (mm_interconnect_0_avalon_spi_max31865_3_s1_address),     //              .address
		.avs_s1_waitrequest (mm_interconnect_0_avalon_spi_max31865_3_s1_waitrequest), //              .waitrequest
		.avs_s1_readdata    (mm_interconnect_0_avalon_spi_max31865_3_s1_readdata),    //              .readdata
		.coe_s2_drdy_n      (avalon_spi_max31865_3_conduit_end_0_drdy_n),             // conduit_end_0.drdy_n
		.coe_s2_sclk        (avalon_spi_max31865_3_conduit_end_0_sclk),               //              .sclk
		.coe_s2_cs_n        (avalon_spi_max31865_3_conduit_end_0_cs_n),               //              .cs_n
		.coe_s2_sdi         (avalon_spi_max31865_3_conduit_end_0_sdi),                //              .sdi
		.coe_s2_sdo         (avalon_spi_max31865_3_conduit_end_0_sdo)                 //              .sdo
	);

	avalon_spi_max31865 #(
		.g_cpol ("'0'")
	) avalon_spi_max31865_4 (
		.csi_clock_clk      (pll_0_sys_clk_clk),                                      //         clock.clk
		.rsi_reset_reset_n  (~rst_controller_reset_out_reset),                        //         reset.reset_n
		.avs_s1_writedata   (mm_interconnect_0_avalon_spi_max31865_4_s1_writedata),   //            s1.writedata
		.avs_s1_read        (mm_interconnect_0_avalon_spi_max31865_4_s1_read),        //              .read
		.avs_s1_write       (mm_interconnect_0_avalon_spi_max31865_4_s1_write),       //              .write
		.avs_s1_address     (mm_interconnect_0_avalon_spi_max31865_4_s1_address),     //              .address
		.avs_s1_waitrequest (mm_interconnect_0_avalon_spi_max31865_4_s1_waitrequest), //              .waitrequest
		.avs_s1_readdata    (mm_interconnect_0_avalon_spi_max31865_4_s1_readdata),    //              .readdata
		.coe_s2_drdy_n      (avalon_spi_max31865_4_conduit_end_0_drdy_n),             // conduit_end_0.drdy_n
		.coe_s2_sclk        (avalon_spi_max31865_4_conduit_end_0_sclk),               //              .sclk
		.coe_s2_cs_n        (avalon_spi_max31865_4_conduit_end_0_cs_n),               //              .cs_n
		.coe_s2_sdi         (avalon_spi_max31865_4_conduit_end_0_sdi),                //              .sdi
		.coe_s2_sdo         (avalon_spi_max31865_4_conduit_end_0_sdo)                 //              .sdo
	);

	avalon_spi_max31865 #(
		.g_cpol ("'0'")
	) avalon_spi_max31865_5 (
		.csi_clock_clk      (pll_0_sys_clk_clk),                                      //         clock.clk
		.rsi_reset_reset_n  (~rst_controller_reset_out_reset),                        //         reset.reset_n
		.avs_s1_writedata   (mm_interconnect_0_avalon_spi_max31865_5_s1_writedata),   //            s1.writedata
		.avs_s1_read        (mm_interconnect_0_avalon_spi_max31865_5_s1_read),        //              .read
		.avs_s1_write       (mm_interconnect_0_avalon_spi_max31865_5_s1_write),       //              .write
		.avs_s1_address     (mm_interconnect_0_avalon_spi_max31865_5_s1_address),     //              .address
		.avs_s1_waitrequest (mm_interconnect_0_avalon_spi_max31865_5_s1_waitrequest), //              .waitrequest
		.avs_s1_readdata    (mm_interconnect_0_avalon_spi_max31865_5_s1_readdata),    //              .readdata
		.coe_s2_drdy_n      (avalon_spi_max31865_5_conduit_end_0_drdy_n),             // conduit_end_0.drdy_n
		.coe_s2_sclk        (avalon_spi_max31865_5_conduit_end_0_sclk),               //              .sclk
		.coe_s2_cs_n        (avalon_spi_max31865_5_conduit_end_0_cs_n),               //              .cs_n
		.coe_s2_sdi         (avalon_spi_max31865_5_conduit_end_0_sdi),                //              .sdi
		.coe_s2_sdo         (avalon_spi_max31865_5_conduit_end_0_sdo)                 //              .sdo
	);

	axi_lw_slave_register #(
		.g_master_id_width   (12),
		.g_master_data_width (32),
		.g_master_addr_width (16)
	) axi_lw_slave_register_0 (
		.rsi_reset_reset_n (~rst_controller_reset_out_reset),                                         //                 reset.reset_n
		.csi_clock_clk     (pll_0_sys_clk_clk),                                                       //                 clock.clk
		.coe_wr_strb       (axi_lw_slave_register_0_conduit_end_0_wr_strb),                           //         conduit_end_0.wr_strb
		.coe_wr_valid      (axi_lw_slave_register_0_conduit_end_0_wr_valid),                          //                      .wr_valid
		.coe_rd_addr       (axi_lw_slave_register_0_conduit_end_0_rd_addr),                           //                      .rd_addr
		.coe_rd_data       (axi_lw_slave_register_0_conduit_end_0_rd_data),                           //                      .rd_data
		.coe_rd_valid      (axi_lw_slave_register_0_conduit_end_0_rd_valid),                          //                      .rd_valid
		.coe_rd_ready      (axi_lw_slave_register_0_conduit_end_0_rd_ready),                          //                      .rd_ready
		.coe_wr_data       (axi_lw_slave_register_0_conduit_end_0_wr_data),                           //                      .wr_data
		.coe_wr_addr       (axi_lw_slave_register_0_conduit_end_0_wr_addr),                           //                      .wr_addr
		.axs_awaddr        (mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_awaddr),  // altera_axi4lite_slave.awaddr
		.axs_awprot        (mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_awprot),  //                      .awprot
		.axs_awvalid       (mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_awvalid), //                      .awvalid
		.axs_awready       (mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_awready), //                      .awready
		.axs_wdata         (mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_wdata),   //                      .wdata
		.axs_wstrb         (mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_wstrb),   //                      .wstrb
		.axs_wvalid        (mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_wvalid),  //                      .wvalid
		.axs_wready        (mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_wready),  //                      .wready
		.axs_bresp         (mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_bresp),   //                      .bresp
		.axs_bvalid        (mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_bvalid),  //                      .bvalid
		.axs_bready        (mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_bready),  //                      .bready
		.axs_araddr        (mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_araddr),  //                      .araddr
		.axs_arprot        (mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_arprot),  //                      .arprot
		.axs_arvalid       (mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_arvalid), //                      .arvalid
		.axs_arready       (mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_arready), //                      .arready
		.axs_rdata         (mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_rdata),   //                      .rdata
		.axs_rresp         (mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_rresp),   //                      .rresp
		.axs_rvalid        (mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_rvalid),  //                      .rvalid
		.axs_rready        (mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_rready)   //                      .rready
	);

	fluid_board_soc_flush_pump_pwm_duty_cycle flush_pump_pwm_duty_cycle (
		.clk        (pll_0_sys_clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                           //               reset.reset_n
		.address    (mm_interconnect_0_flush_pump_pwm_duty_cycle_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_flush_pump_pwm_duty_cycle_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_flush_pump_pwm_duty_cycle_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_flush_pump_pwm_duty_cycle_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_flush_pump_pwm_duty_cycle_s1_readdata),   //                    .readdata
		.out_port   (flush_pump_pwm_duty_cycle_external_connection_export)       // external_connection.export
	);

	fluid_board_soc_flush_pump_pwm_duty_cycle flush_pump_pwm_freq (
		.clk        (pll_0_sys_clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                     //               reset.reset_n
		.address    (mm_interconnect_0_flush_pump_pwm_freq_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_flush_pump_pwm_freq_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_flush_pump_pwm_freq_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_flush_pump_pwm_freq_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_flush_pump_pwm_freq_s1_readdata),   //                    .readdata
		.out_port   (flush_pump_pwm_freq_external_connection_export)       // external_connection.export
	);

	fluid_board_soc_fpga_only_master #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) fpga_only_master (
		.clk_clk              (pll_0_sys_clk_clk),                     //          clk.clk
		.clk_reset_reset      (~qsys_reset_reset_n),                   //    clk_reset.reset
		.master_address       (fpga_only_master_master_address),       //       master.address
		.master_readdata      (fpga_only_master_master_readdata),      //             .readdata
		.master_read          (fpga_only_master_master_read),          //             .read
		.master_write         (fpga_only_master_master_write),         //             .write
		.master_writedata     (fpga_only_master_master_writedata),     //             .writedata
		.master_waitrequest   (fpga_only_master_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (fpga_only_master_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (fpga_only_master_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                                       // master_reset.reset
	);

	fluid_board_soc_hps_0 #(
		.F2S_Width (0),
		.S2F_Width (2)
	) hps_0 (
		.uart1_cts                (hps_0_uart1_cts),                 //             uart1.cts
		.uart1_dsr                (hps_0_uart1_dsr),                 //                  .dsr
		.uart1_dcd                (hps_0_uart1_dcd),                 //                  .dcd
		.uart1_ri                 (hps_0_uart1_ri),                  //                  .ri
		.uart1_dtr                (hps_0_uart1_dtr),                 //                  .dtr
		.uart1_rts                (hps_0_uart1_rts),                 //                  .rts
		.uart1_out1_n             (hps_0_uart1_out1_n),              //                  .out1_n
		.uart1_out2_n             (hps_0_uart1_out2_n),              //                  .out2_n
		.uart1_rxd                (hps_0_uart1_rxd),                 //                  .rxd
		.uart1_txd                (hps_0_uart1_txd),                 //                  .txd
		.mem_a                    (memory_mem_a),                    //            memory.mem_a
		.mem_ba                   (memory_mem_ba),                   //                  .mem_ba
		.mem_ck                   (memory_mem_ck),                   //                  .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),                 //                  .mem_ck_n
		.mem_cke                  (memory_mem_cke),                  //                  .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),                 //                  .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),                //                  .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),                //                  .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),                 //                  .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),              //                  .mem_reset_n
		.mem_dq                   (memory_mem_dq),                   //                  .mem_dq
		.mem_dqs                  (memory_mem_dqs),                  //                  .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),                //                  .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                  //                  .mem_odt
		.mem_dm                   (memory_mem_dm),                   //                  .mem_dm
		.oct_rzqin                (memory_oct_rzqin),                //                  .oct_rzqin
		.hps_io_emac0_inst_TX_CLK (hps_io_hps_io_emac0_inst_TX_CLK), //            hps_io.hps_io_emac0_inst_TX_CLK
		.hps_io_emac0_inst_TXD0   (hps_io_hps_io_emac0_inst_TXD0),   //                  .hps_io_emac0_inst_TXD0
		.hps_io_emac0_inst_TXD1   (hps_io_hps_io_emac0_inst_TXD1),   //                  .hps_io_emac0_inst_TXD1
		.hps_io_emac0_inst_TXD2   (hps_io_hps_io_emac0_inst_TXD2),   //                  .hps_io_emac0_inst_TXD2
		.hps_io_emac0_inst_TXD3   (hps_io_hps_io_emac0_inst_TXD3),   //                  .hps_io_emac0_inst_TXD3
		.hps_io_emac0_inst_RXD0   (hps_io_hps_io_emac0_inst_RXD0),   //                  .hps_io_emac0_inst_RXD0
		.hps_io_emac0_inst_MDIO   (hps_io_hps_io_emac0_inst_MDIO),   //                  .hps_io_emac0_inst_MDIO
		.hps_io_emac0_inst_MDC    (hps_io_hps_io_emac0_inst_MDC),    //                  .hps_io_emac0_inst_MDC
		.hps_io_emac0_inst_RX_CTL (hps_io_hps_io_emac0_inst_RX_CTL), //                  .hps_io_emac0_inst_RX_CTL
		.hps_io_emac0_inst_TX_CTL (hps_io_hps_io_emac0_inst_TX_CTL), //                  .hps_io_emac0_inst_TX_CTL
		.hps_io_emac0_inst_RX_CLK (hps_io_hps_io_emac0_inst_RX_CLK), //                  .hps_io_emac0_inst_RX_CLK
		.hps_io_emac0_inst_RXD1   (hps_io_hps_io_emac0_inst_RXD1),   //                  .hps_io_emac0_inst_RXD1
		.hps_io_emac0_inst_RXD2   (hps_io_hps_io_emac0_inst_RXD2),   //                  .hps_io_emac0_inst_RXD2
		.hps_io_emac0_inst_RXD3   (hps_io_hps_io_emac0_inst_RXD3),   //                  .hps_io_emac0_inst_RXD3
		.hps_io_sdio_inst_CMD     (hps_io_hps_io_sdio_inst_CMD),     //                  .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_io_hps_io_sdio_inst_D0),      //                  .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_io_hps_io_sdio_inst_D1),      //                  .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_D4      (hps_io_hps_io_sdio_inst_D4),      //                  .hps_io_sdio_inst_D4
		.hps_io_sdio_inst_D5      (hps_io_hps_io_sdio_inst_D5),      //                  .hps_io_sdio_inst_D5
		.hps_io_sdio_inst_D6      (hps_io_hps_io_sdio_inst_D6),      //                  .hps_io_sdio_inst_D6
		.hps_io_sdio_inst_D7      (hps_io_hps_io_sdio_inst_D7),      //                  .hps_io_sdio_inst_D7
		.hps_io_sdio_inst_CLK     (hps_io_hps_io_sdio_inst_CLK),     //                  .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_io_hps_io_sdio_inst_D2),      //                  .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_io_hps_io_sdio_inst_D3),      //                  .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_io_hps_io_usb1_inst_D0),      //                  .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_io_hps_io_usb1_inst_D1),      //                  .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_io_hps_io_usb1_inst_D2),      //                  .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_io_hps_io_usb1_inst_D3),      //                  .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_io_hps_io_usb1_inst_D4),      //                  .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_io_hps_io_usb1_inst_D5),      //                  .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_io_hps_io_usb1_inst_D6),      //                  .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_io_hps_io_usb1_inst_D7),      //                  .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_io_hps_io_usb1_inst_CLK),     //                  .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_io_hps_io_usb1_inst_STP),     //                  .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_io_hps_io_usb1_inst_DIR),     //                  .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_io_hps_io_usb1_inst_NXT),     //                  .hps_io_usb1_inst_NXT
		.hps_io_uart0_inst_RX     (hps_io_hps_io_uart0_inst_RX),     //                  .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_io_hps_io_uart0_inst_TX),     //                  .hps_io_uart0_inst_TX
		.hps_io_gpio_inst_GPIO37  (hps_io_hps_io_gpio_inst_GPIO37),  //                  .hps_io_gpio_inst_GPIO37
		.hps_io_gpio_inst_GPIO44  (hps_io_hps_io_gpio_inst_GPIO44),  //                  .hps_io_gpio_inst_GPIO44
		.hps_io_gpio_inst_GPIO59  (hps_io_hps_io_gpio_inst_GPIO59),  //                  .hps_io_gpio_inst_GPIO59
		.h2f_rst_n                (hps_0_h2f_reset_reset),           //         h2f_reset.reset_n
		.h2f_axi_clk              (pll_0_sys_clk_clk),               //     h2f_axi_clock.clk
		.h2f_AWID                 (hps_0_h2f_axi_master_awid),       //    h2f_axi_master.awid
		.h2f_AWADDR               (hps_0_h2f_axi_master_awaddr),     //                  .awaddr
		.h2f_AWLEN                (hps_0_h2f_axi_master_awlen),      //                  .awlen
		.h2f_AWSIZE               (hps_0_h2f_axi_master_awsize),     //                  .awsize
		.h2f_AWBURST              (hps_0_h2f_axi_master_awburst),    //                  .awburst
		.h2f_AWLOCK               (hps_0_h2f_axi_master_awlock),     //                  .awlock
		.h2f_AWCACHE              (hps_0_h2f_axi_master_awcache),    //                  .awcache
		.h2f_AWPROT               (hps_0_h2f_axi_master_awprot),     //                  .awprot
		.h2f_AWVALID              (hps_0_h2f_axi_master_awvalid),    //                  .awvalid
		.h2f_AWREADY              (hps_0_h2f_axi_master_awready),    //                  .awready
		.h2f_WID                  (hps_0_h2f_axi_master_wid),        //                  .wid
		.h2f_WDATA                (hps_0_h2f_axi_master_wdata),      //                  .wdata
		.h2f_WSTRB                (hps_0_h2f_axi_master_wstrb),      //                  .wstrb
		.h2f_WLAST                (hps_0_h2f_axi_master_wlast),      //                  .wlast
		.h2f_WVALID               (hps_0_h2f_axi_master_wvalid),     //                  .wvalid
		.h2f_WREADY               (hps_0_h2f_axi_master_wready),     //                  .wready
		.h2f_BID                  (hps_0_h2f_axi_master_bid),        //                  .bid
		.h2f_BRESP                (hps_0_h2f_axi_master_bresp),      //                  .bresp
		.h2f_BVALID               (hps_0_h2f_axi_master_bvalid),     //                  .bvalid
		.h2f_BREADY               (hps_0_h2f_axi_master_bready),     //                  .bready
		.h2f_ARID                 (hps_0_h2f_axi_master_arid),       //                  .arid
		.h2f_ARADDR               (hps_0_h2f_axi_master_araddr),     //                  .araddr
		.h2f_ARLEN                (hps_0_h2f_axi_master_arlen),      //                  .arlen
		.h2f_ARSIZE               (hps_0_h2f_axi_master_arsize),     //                  .arsize
		.h2f_ARBURST              (hps_0_h2f_axi_master_arburst),    //                  .arburst
		.h2f_ARLOCK               (hps_0_h2f_axi_master_arlock),     //                  .arlock
		.h2f_ARCACHE              (hps_0_h2f_axi_master_arcache),    //                  .arcache
		.h2f_ARPROT               (hps_0_h2f_axi_master_arprot),     //                  .arprot
		.h2f_ARVALID              (hps_0_h2f_axi_master_arvalid),    //                  .arvalid
		.h2f_ARREADY              (hps_0_h2f_axi_master_arready),    //                  .arready
		.h2f_RID                  (hps_0_h2f_axi_master_rid),        //                  .rid
		.h2f_RDATA                (hps_0_h2f_axi_master_rdata),      //                  .rdata
		.h2f_RRESP                (hps_0_h2f_axi_master_rresp),      //                  .rresp
		.h2f_RLAST                (hps_0_h2f_axi_master_rlast),      //                  .rlast
		.h2f_RVALID               (hps_0_h2f_axi_master_rvalid),     //                  .rvalid
		.h2f_RREADY               (hps_0_h2f_axi_master_rready),     //                  .rready
		.h2f_lw_axi_clk           (pll_0_sys_clk_clk),               //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (hps_0_h2f_lw_axi_master_awid),    // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (hps_0_h2f_lw_axi_master_awaddr),  //                  .awaddr
		.h2f_lw_AWLEN             (hps_0_h2f_lw_axi_master_awlen),   //                  .awlen
		.h2f_lw_AWSIZE            (hps_0_h2f_lw_axi_master_awsize),  //                  .awsize
		.h2f_lw_AWBURST           (hps_0_h2f_lw_axi_master_awburst), //                  .awburst
		.h2f_lw_AWLOCK            (hps_0_h2f_lw_axi_master_awlock),  //                  .awlock
		.h2f_lw_AWCACHE           (hps_0_h2f_lw_axi_master_awcache), //                  .awcache
		.h2f_lw_AWPROT            (hps_0_h2f_lw_axi_master_awprot),  //                  .awprot
		.h2f_lw_AWVALID           (hps_0_h2f_lw_axi_master_awvalid), //                  .awvalid
		.h2f_lw_AWREADY           (hps_0_h2f_lw_axi_master_awready), //                  .awready
		.h2f_lw_WID               (hps_0_h2f_lw_axi_master_wid),     //                  .wid
		.h2f_lw_WDATA             (hps_0_h2f_lw_axi_master_wdata),   //                  .wdata
		.h2f_lw_WSTRB             (hps_0_h2f_lw_axi_master_wstrb),   //                  .wstrb
		.h2f_lw_WLAST             (hps_0_h2f_lw_axi_master_wlast),   //                  .wlast
		.h2f_lw_WVALID            (hps_0_h2f_lw_axi_master_wvalid),  //                  .wvalid
		.h2f_lw_WREADY            (hps_0_h2f_lw_axi_master_wready),  //                  .wready
		.h2f_lw_BID               (hps_0_h2f_lw_axi_master_bid),     //                  .bid
		.h2f_lw_BRESP             (hps_0_h2f_lw_axi_master_bresp),   //                  .bresp
		.h2f_lw_BVALID            (hps_0_h2f_lw_axi_master_bvalid),  //                  .bvalid
		.h2f_lw_BREADY            (hps_0_h2f_lw_axi_master_bready),  //                  .bready
		.h2f_lw_ARID              (hps_0_h2f_lw_axi_master_arid),    //                  .arid
		.h2f_lw_ARADDR            (hps_0_h2f_lw_axi_master_araddr),  //                  .araddr
		.h2f_lw_ARLEN             (hps_0_h2f_lw_axi_master_arlen),   //                  .arlen
		.h2f_lw_ARSIZE            (hps_0_h2f_lw_axi_master_arsize),  //                  .arsize
		.h2f_lw_ARBURST           (hps_0_h2f_lw_axi_master_arburst), //                  .arburst
		.h2f_lw_ARLOCK            (hps_0_h2f_lw_axi_master_arlock),  //                  .arlock
		.h2f_lw_ARCACHE           (hps_0_h2f_lw_axi_master_arcache), //                  .arcache
		.h2f_lw_ARPROT            (hps_0_h2f_lw_axi_master_arprot),  //                  .arprot
		.h2f_lw_ARVALID           (hps_0_h2f_lw_axi_master_arvalid), //                  .arvalid
		.h2f_lw_ARREADY           (hps_0_h2f_lw_axi_master_arready), //                  .arready
		.h2f_lw_RID               (hps_0_h2f_lw_axi_master_rid),     //                  .rid
		.h2f_lw_RDATA             (hps_0_h2f_lw_axi_master_rdata),   //                  .rdata
		.h2f_lw_RRESP             (hps_0_h2f_lw_axi_master_rresp),   //                  .rresp
		.h2f_lw_RLAST             (hps_0_h2f_lw_axi_master_rlast),   //                  .rlast
		.h2f_lw_RVALID            (hps_0_h2f_lw_axi_master_rvalid),  //                  .rvalid
		.h2f_lw_RREADY            (hps_0_h2f_lw_axi_master_rready),  //                  .rready
		.f2h_irq_p0               (hps_0_f2h_irq0_irq),              //          f2h_irq0.irq
		.f2h_irq_p1               (hps_0_f2h_irq1_irq)               //          f2h_irq1.irq
	);

	i2c_opencores i2c_master_d (
		.sda_pad_io (i2c_master_d_conduit_end_sda),                            //      conduit_end.sda
		.scl_pad_io (i2c_master_d_conduit_end_scl),                            //                 .scl
		.wb_inta_o  (irq_mapper_002_receiver6_irq),                            // interrupt_sender.irq
		.wb_dat_o   (mm_interconnect_0_i2c_master_d_avalon_slave_readdata),    //     avalon_slave.readdata
		.wb_stb_i   (mm_interconnect_0_i2c_master_d_avalon_slave_chipselect),  //                 .chipselect
		.wb_ack_o   (mm_interconnect_0_i2c_master_d_avalon_slave_waitrequest), //                 .waitrequest_n
		.wb_adr_i   (mm_interconnect_0_i2c_master_d_avalon_slave_address),     //                 .address
		.wb_we_i    (mm_interconnect_0_i2c_master_d_avalon_slave_write),       //                 .write
		.wb_dat_i   (mm_interconnect_0_i2c_master_d_avalon_slave_writedata),   //                 .writedata
		.wb_clk_i   (pll_0_sys_clk_clk),                                       //            clock.clk
		.wb_rst_i   (rst_controller_reset_out_reset)                           //      clock_reset.reset
	);

	i2c_opencores i2c_master_f (
		.sda_pad_io (i2c_master_f_conduit_end_sda),                            //      conduit_end.sda
		.scl_pad_io (i2c_master_f_conduit_end_scl),                            //                 .scl
		.wb_inta_o  (irq_mapper_002_receiver5_irq),                            // interrupt_sender.irq
		.wb_dat_o   (mm_interconnect_0_i2c_master_f_avalon_slave_readdata),    //     avalon_slave.readdata
		.wb_stb_i   (mm_interconnect_0_i2c_master_f_avalon_slave_chipselect),  //                 .chipselect
		.wb_ack_o   (mm_interconnect_0_i2c_master_f_avalon_slave_waitrequest), //                 .waitrequest_n
		.wb_adr_i   (mm_interconnect_0_i2c_master_f_avalon_slave_address),     //                 .address
		.wb_we_i    (mm_interconnect_0_i2c_master_f_avalon_slave_write),       //                 .write
		.wb_dat_i   (mm_interconnect_0_i2c_master_f_avalon_slave_writedata),   //                 .writedata
		.wb_clk_i   (pll_0_sys_clk_clk),                                       //            clock.clk
		.wb_rst_i   (rst_controller_reset_out_reset)                           //      clock_reset.reset
	);

	i2c_opencores i2c_master_is1 (
		.sda_pad_io (i2c_master_is1_conduit_end_sda),                            //      conduit_end.sda
		.scl_pad_io (i2c_master_is1_conduit_end_scl),                            //                 .scl
		.wb_inta_o  (irq_mapper_002_receiver0_irq),                              // interrupt_sender.irq
		.wb_dat_o   (mm_interconnect_0_i2c_master_is1_avalon_slave_readdata),    //     avalon_slave.readdata
		.wb_stb_i   (mm_interconnect_0_i2c_master_is1_avalon_slave_chipselect),  //                 .chipselect
		.wb_ack_o   (mm_interconnect_0_i2c_master_is1_avalon_slave_waitrequest), //                 .waitrequest_n
		.wb_adr_i   (mm_interconnect_0_i2c_master_is1_avalon_slave_address),     //                 .address
		.wb_we_i    (mm_interconnect_0_i2c_master_is1_avalon_slave_write),       //                 .write
		.wb_dat_i   (mm_interconnect_0_i2c_master_is1_avalon_slave_writedata),   //                 .writedata
		.wb_clk_i   (pll_0_sys_clk_clk),                                         //            clock.clk
		.wb_rst_i   (rst_controller_reset_out_reset)                             //      clock_reset.reset
	);

	i2c_opencores i2c_master_is2 (
		.sda_pad_io (i2c_master_is2_conduit_end_sda),                            //      conduit_end.sda
		.scl_pad_io (i2c_master_is2_conduit_end_scl),                            //                 .scl
		.wb_inta_o  (irq_mapper_002_receiver1_irq),                              // interrupt_sender.irq
		.wb_dat_o   (mm_interconnect_0_i2c_master_is2_avalon_slave_readdata),    //     avalon_slave.readdata
		.wb_stb_i   (mm_interconnect_0_i2c_master_is2_avalon_slave_chipselect),  //                 .chipselect
		.wb_ack_o   (mm_interconnect_0_i2c_master_is2_avalon_slave_waitrequest), //                 .waitrequest_n
		.wb_adr_i   (mm_interconnect_0_i2c_master_is2_avalon_slave_address),     //                 .address
		.wb_we_i    (mm_interconnect_0_i2c_master_is2_avalon_slave_write),       //                 .write
		.wb_dat_i   (mm_interconnect_0_i2c_master_is2_avalon_slave_writedata),   //                 .writedata
		.wb_clk_i   (pll_0_sys_clk_clk),                                         //            clock.clk
		.wb_rst_i   (rst_controller_reset_out_reset)                             //      clock_reset.reset
	);

	i2c_opencores i2c_master_is3 (
		.sda_pad_io (i2c_master_is3_conduit_end_sda),                            //      conduit_end.sda
		.scl_pad_io (i2c_master_is3_conduit_end_scl),                            //                 .scl
		.wb_inta_o  (irq_mapper_002_receiver2_irq),                              // interrupt_sender.irq
		.wb_dat_o   (mm_interconnect_0_i2c_master_is3_avalon_slave_readdata),    //     avalon_slave.readdata
		.wb_stb_i   (mm_interconnect_0_i2c_master_is3_avalon_slave_chipselect),  //                 .chipselect
		.wb_ack_o   (mm_interconnect_0_i2c_master_is3_avalon_slave_waitrequest), //                 .waitrequest_n
		.wb_adr_i   (mm_interconnect_0_i2c_master_is3_avalon_slave_address),     //                 .address
		.wb_we_i    (mm_interconnect_0_i2c_master_is3_avalon_slave_write),       //                 .write
		.wb_dat_i   (mm_interconnect_0_i2c_master_is3_avalon_slave_writedata),   //                 .writedata
		.wb_clk_i   (pll_0_sys_clk_clk),                                         //            clock.clk
		.wb_rst_i   (rst_controller_reset_out_reset)                             //      clock_reset.reset
	);

	i2c_opencores i2c_master_is4 (
		.sda_pad_io (i2c_master_is4_conduit_end_sda),                            //      conduit_end.sda
		.scl_pad_io (i2c_master_is4_conduit_end_scl),                            //                 .scl
		.wb_inta_o  (irq_mapper_002_receiver3_irq),                              // interrupt_sender.irq
		.wb_dat_o   (mm_interconnect_0_i2c_master_is4_avalon_slave_readdata),    //     avalon_slave.readdata
		.wb_stb_i   (mm_interconnect_0_i2c_master_is4_avalon_slave_chipselect),  //                 .chipselect
		.wb_ack_o   (mm_interconnect_0_i2c_master_is4_avalon_slave_waitrequest), //                 .waitrequest_n
		.wb_adr_i   (mm_interconnect_0_i2c_master_is4_avalon_slave_address),     //                 .address
		.wb_we_i    (mm_interconnect_0_i2c_master_is4_avalon_slave_write),       //                 .write
		.wb_dat_i   (mm_interconnect_0_i2c_master_is4_avalon_slave_writedata),   //                 .writedata
		.wb_clk_i   (pll_0_sys_clk_clk),                                         //            clock.clk
		.wb_rst_i   (rst_controller_reset_out_reset)                             //      clock_reset.reset
	);

	i2c_opencores i2c_master_p (
		.sda_pad_io (i2c_master_p_conduit_end_sda),                            //      conduit_end.sda
		.scl_pad_io (i2c_master_p_conduit_end_scl),                            //                 .scl
		.wb_inta_o  (irq_mapper_002_receiver4_irq),                            // interrupt_sender.irq
		.wb_dat_o   (mm_interconnect_0_i2c_master_p_avalon_slave_readdata),    //     avalon_slave.readdata
		.wb_stb_i   (mm_interconnect_0_i2c_master_p_avalon_slave_chipselect),  //                 .chipselect
		.wb_ack_o   (mm_interconnect_0_i2c_master_p_avalon_slave_waitrequest), //                 .waitrequest_n
		.wb_adr_i   (mm_interconnect_0_i2c_master_p_avalon_slave_address),     //                 .address
		.wb_we_i    (mm_interconnect_0_i2c_master_p_avalon_slave_write),       //                 .write
		.wb_dat_i   (mm_interconnect_0_i2c_master_p_avalon_slave_writedata),   //                 .writedata
		.wb_clk_i   (pll_0_sys_clk_clk),                                       //            clock.clk
		.wb_rst_i   (rst_controller_reset_out_reset)                           //      clock_reset.reset
	);

	fluid_board_soc_jtag_uart jtag_uart (
		.clk            (pll_0_sys_clk_clk),                                         //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	fluid_board_soc_nios2_qsys_0 nios2_qsys_0 (
		.clk                                 (pll_0_sys_clk_clk),                                          //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_qsys_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_qsys_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_qsys_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_qsys_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_qsys_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_qsys_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_qsys_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_qsys_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_qsys_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_qsys_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_qsys_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_qsys_0_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_qsys_0_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_qsys_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                           //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       (),                                                           // custom_instruction_master.readra
		.cpu_resetrequest                    (nios2_qsys_0_cpu_resetrequest_conduit_cpu_resetrequest),     //  cpu_resetrequest_conduit.cpu_resetrequest
		.cpu_resettaken                      (nios2_qsys_0_cpu_resetrequest_conduit_cpu_resettaken)        //                          .cpu_resettaken
	);

	fluid_board_soc_onchip_memory_nios_arm onchip_memory_nios_arm (
		.address     (mm_interconnect_0_onchip_memory_nios_arm_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_onchip_memory_nios_arm_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_onchip_memory_nios_arm_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_onchip_memory_nios_arm_s1_write),      //       .write
		.readdata    (mm_interconnect_0_onchip_memory_nios_arm_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_onchip_memory_nios_arm_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_onchip_memory_nios_arm_s1_byteenable), //       .byteenable
		.address2    (mm_interconnect_0_onchip_memory_nios_arm_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_onchip_memory_nios_arm_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_onchip_memory_nios_arm_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_onchip_memory_nios_arm_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_onchip_memory_nios_arm_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_onchip_memory_nios_arm_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_onchip_memory_nios_arm_s2_byteenable), //       .byteenable
		.clk         (pll_0_sys_clk_clk),                                      //   clk1.clk
		.reset       (rst_controller_001_reset_out_reset),                     // reset1.reset
		.reset_req   (rst_controller_001_reset_out_reset_req)                  //       .reset_req
	);

	fluid_board_soc_onchip_memory_nios_cpu onchip_memory_nios_cpu (
		.address     (mm_interconnect_0_onchip_memory_nios_cpu_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_onchip_memory_nios_cpu_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_onchip_memory_nios_cpu_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_onchip_memory_nios_cpu_s1_write),      //       .write
		.readdata    (mm_interconnect_0_onchip_memory_nios_cpu_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_onchip_memory_nios_cpu_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_onchip_memory_nios_cpu_s1_byteenable), //       .byteenable
		.address2    (mm_interconnect_0_onchip_memory_nios_cpu_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_onchip_memory_nios_cpu_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_onchip_memory_nios_cpu_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_onchip_memory_nios_cpu_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_onchip_memory_nios_cpu_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_onchip_memory_nios_cpu_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_onchip_memory_nios_cpu_s2_byteenable), //       .byteenable
		.clk         (pll_0_sys_clk_clk),                                      //   clk1.clk
		.reset       (rst_controller_001_reset_out_reset),                     // reset1.reset
		.reset_req   (rst_controller_001_reset_out_reset_req)                  //       .reset_req
	);

	fluid_board_soc_pio_input pio_input (
		.clk        (pll_0_sys_clk_clk),                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_pio_input_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_input_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_input_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_input_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_input_s1_readdata),   //                    .readdata
		.in_port    (pio_input_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_002_receiver9_irq)               //                 irq.irq
	);

	fluid_board_soc_pio_output pio_output (
		.clk        (pll_0_sys_clk_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_pio_output_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_output_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_output_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_output_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_output_s1_readdata),   //                    .readdata
		.out_port   (pio_output_external_connection_export)       // external_connection.export
	);

	fluid_board_soc_pio_reset_nios pio_reset_nios (
		.clk        (pll_0_sys_clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_pio_reset_nios_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_reset_nios_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_reset_nios_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_reset_nios_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_reset_nios_s1_readdata),   //                    .readdata
		.out_port   (pio_reset_nios_external_connection_export)       // external_connection.export
	);

	fluid_board_soc_flush_pump_pwm_duty_cycle pio_watchdog_cnt (
		.clk        (pll_0_sys_clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_0_pio_watchdog_cnt_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_watchdog_cnt_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_watchdog_cnt_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_watchdog_cnt_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_watchdog_cnt_s1_readdata),   //                    .readdata
		.out_port   (pio_watchdog_cnt_external_connection_export)       // external_connection.export
	);

	fluid_board_soc_flush_pump_pwm_duty_cycle pio_watchdog_freq (
		.clk        (pll_0_sys_clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (mm_interconnect_0_pio_watchdog_freq_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_watchdog_freq_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_watchdog_freq_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_watchdog_freq_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_watchdog_freq_s1_readdata),   //                    .readdata
		.out_port   (pio_watchdog_freq_external_connection_export)       // external_connection.export
	);

	fluid_board_soc_pll_0 pll_0 (
		.refclk   (pll_0_refclk_clk),    //  refclk.clk
		.rst      (pll_0_reset_reset),   //   reset.reset
		.outclk_0 (pll_0_sys_clk_clk),   // outclk0.clk
		.locked   (pll_0_locked_export)  //  locked.export
	);

	fluid_board_soc_sysid sysid (
		.clock    (pll_0_sys_clk_clk),                              //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),            //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	fluid_board_soc_timer_0 timer_0 (
		.clk        (pll_0_sys_clk_clk),                       //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_002_receiver7_irq)             //   irq.irq
	);

	fluid_board_soc_timer_0 timer_1 (
		.clk        (pll_0_sys_clk_clk),                       //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_1_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_1_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_1_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_1_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_1_s1_write),     //      .write_n
		.irq        (irq_mapper_002_receiver8_irq)             //   irq.irq
	);

	fluid_board_soc_timer_0 timer_2 (
		.clk        (pll_0_sys_clk_clk),                       //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_2_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_2_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_2_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_2_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_2_s1_write),     //      .write_n
		.irq        (irq_mapper_002_receiver11_irq)            //   irq.irq
	);

	fluid_board_soc_mm_interconnect_0 mm_interconnect_0 (
		.axi_lw_slave_register_0_altera_axi4lite_slave_awaddr             (mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_awaddr),  //              axi_lw_slave_register_0_altera_axi4lite_slave.awaddr
		.axi_lw_slave_register_0_altera_axi4lite_slave_awprot             (mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_awprot),  //                                                           .awprot
		.axi_lw_slave_register_0_altera_axi4lite_slave_awvalid            (mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_awvalid), //                                                           .awvalid
		.axi_lw_slave_register_0_altera_axi4lite_slave_awready            (mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_awready), //                                                           .awready
		.axi_lw_slave_register_0_altera_axi4lite_slave_wdata              (mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_wdata),   //                                                           .wdata
		.axi_lw_slave_register_0_altera_axi4lite_slave_wstrb              (mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_wstrb),   //                                                           .wstrb
		.axi_lw_slave_register_0_altera_axi4lite_slave_wvalid             (mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_wvalid),  //                                                           .wvalid
		.axi_lw_slave_register_0_altera_axi4lite_slave_wready             (mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_wready),  //                                                           .wready
		.axi_lw_slave_register_0_altera_axi4lite_slave_bresp              (mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_bresp),   //                                                           .bresp
		.axi_lw_slave_register_0_altera_axi4lite_slave_bvalid             (mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_bvalid),  //                                                           .bvalid
		.axi_lw_slave_register_0_altera_axi4lite_slave_bready             (mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_bready),  //                                                           .bready
		.axi_lw_slave_register_0_altera_axi4lite_slave_araddr             (mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_araddr),  //                                                           .araddr
		.axi_lw_slave_register_0_altera_axi4lite_slave_arprot             (mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_arprot),  //                                                           .arprot
		.axi_lw_slave_register_0_altera_axi4lite_slave_arvalid            (mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_arvalid), //                                                           .arvalid
		.axi_lw_slave_register_0_altera_axi4lite_slave_arready            (mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_arready), //                                                           .arready
		.axi_lw_slave_register_0_altera_axi4lite_slave_rdata              (mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_rdata),   //                                                           .rdata
		.axi_lw_slave_register_0_altera_axi4lite_slave_rresp              (mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_rresp),   //                                                           .rresp
		.axi_lw_slave_register_0_altera_axi4lite_slave_rvalid             (mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_rvalid),  //                                                           .rvalid
		.axi_lw_slave_register_0_altera_axi4lite_slave_rready             (mm_interconnect_0_axi_lw_slave_register_0_altera_axi4lite_slave_rready),  //                                                           .rready
		.hps_0_h2f_axi_master_awid                                        (hps_0_h2f_axi_master_awid),                                               //                                       hps_0_h2f_axi_master.awid
		.hps_0_h2f_axi_master_awaddr                                      (hps_0_h2f_axi_master_awaddr),                                             //                                                           .awaddr
		.hps_0_h2f_axi_master_awlen                                       (hps_0_h2f_axi_master_awlen),                                              //                                                           .awlen
		.hps_0_h2f_axi_master_awsize                                      (hps_0_h2f_axi_master_awsize),                                             //                                                           .awsize
		.hps_0_h2f_axi_master_awburst                                     (hps_0_h2f_axi_master_awburst),                                            //                                                           .awburst
		.hps_0_h2f_axi_master_awlock                                      (hps_0_h2f_axi_master_awlock),                                             //                                                           .awlock
		.hps_0_h2f_axi_master_awcache                                     (hps_0_h2f_axi_master_awcache),                                            //                                                           .awcache
		.hps_0_h2f_axi_master_awprot                                      (hps_0_h2f_axi_master_awprot),                                             //                                                           .awprot
		.hps_0_h2f_axi_master_awvalid                                     (hps_0_h2f_axi_master_awvalid),                                            //                                                           .awvalid
		.hps_0_h2f_axi_master_awready                                     (hps_0_h2f_axi_master_awready),                                            //                                                           .awready
		.hps_0_h2f_axi_master_wid                                         (hps_0_h2f_axi_master_wid),                                                //                                                           .wid
		.hps_0_h2f_axi_master_wdata                                       (hps_0_h2f_axi_master_wdata),                                              //                                                           .wdata
		.hps_0_h2f_axi_master_wstrb                                       (hps_0_h2f_axi_master_wstrb),                                              //                                                           .wstrb
		.hps_0_h2f_axi_master_wlast                                       (hps_0_h2f_axi_master_wlast),                                              //                                                           .wlast
		.hps_0_h2f_axi_master_wvalid                                      (hps_0_h2f_axi_master_wvalid),                                             //                                                           .wvalid
		.hps_0_h2f_axi_master_wready                                      (hps_0_h2f_axi_master_wready),                                             //                                                           .wready
		.hps_0_h2f_axi_master_bid                                         (hps_0_h2f_axi_master_bid),                                                //                                                           .bid
		.hps_0_h2f_axi_master_bresp                                       (hps_0_h2f_axi_master_bresp),                                              //                                                           .bresp
		.hps_0_h2f_axi_master_bvalid                                      (hps_0_h2f_axi_master_bvalid),                                             //                                                           .bvalid
		.hps_0_h2f_axi_master_bready                                      (hps_0_h2f_axi_master_bready),                                             //                                                           .bready
		.hps_0_h2f_axi_master_arid                                        (hps_0_h2f_axi_master_arid),                                               //                                                           .arid
		.hps_0_h2f_axi_master_araddr                                      (hps_0_h2f_axi_master_araddr),                                             //                                                           .araddr
		.hps_0_h2f_axi_master_arlen                                       (hps_0_h2f_axi_master_arlen),                                              //                                                           .arlen
		.hps_0_h2f_axi_master_arsize                                      (hps_0_h2f_axi_master_arsize),                                             //                                                           .arsize
		.hps_0_h2f_axi_master_arburst                                     (hps_0_h2f_axi_master_arburst),                                            //                                                           .arburst
		.hps_0_h2f_axi_master_arlock                                      (hps_0_h2f_axi_master_arlock),                                             //                                                           .arlock
		.hps_0_h2f_axi_master_arcache                                     (hps_0_h2f_axi_master_arcache),                                            //                                                           .arcache
		.hps_0_h2f_axi_master_arprot                                      (hps_0_h2f_axi_master_arprot),                                             //                                                           .arprot
		.hps_0_h2f_axi_master_arvalid                                     (hps_0_h2f_axi_master_arvalid),                                            //                                                           .arvalid
		.hps_0_h2f_axi_master_arready                                     (hps_0_h2f_axi_master_arready),                                            //                                                           .arready
		.hps_0_h2f_axi_master_rid                                         (hps_0_h2f_axi_master_rid),                                                //                                                           .rid
		.hps_0_h2f_axi_master_rdata                                       (hps_0_h2f_axi_master_rdata),                                              //                                                           .rdata
		.hps_0_h2f_axi_master_rresp                                       (hps_0_h2f_axi_master_rresp),                                              //                                                           .rresp
		.hps_0_h2f_axi_master_rlast                                       (hps_0_h2f_axi_master_rlast),                                              //                                                           .rlast
		.hps_0_h2f_axi_master_rvalid                                      (hps_0_h2f_axi_master_rvalid),                                             //                                                           .rvalid
		.hps_0_h2f_axi_master_rready                                      (hps_0_h2f_axi_master_rready),                                             //                                                           .rready
		.hps_0_h2f_lw_axi_master_awid                                     (hps_0_h2f_lw_axi_master_awid),                                            //                                    hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                                   (hps_0_h2f_lw_axi_master_awaddr),                                          //                                                           .awaddr
		.hps_0_h2f_lw_axi_master_awlen                                    (hps_0_h2f_lw_axi_master_awlen),                                           //                                                           .awlen
		.hps_0_h2f_lw_axi_master_awsize                                   (hps_0_h2f_lw_axi_master_awsize),                                          //                                                           .awsize
		.hps_0_h2f_lw_axi_master_awburst                                  (hps_0_h2f_lw_axi_master_awburst),                                         //                                                           .awburst
		.hps_0_h2f_lw_axi_master_awlock                                   (hps_0_h2f_lw_axi_master_awlock),                                          //                                                           .awlock
		.hps_0_h2f_lw_axi_master_awcache                                  (hps_0_h2f_lw_axi_master_awcache),                                         //                                                           .awcache
		.hps_0_h2f_lw_axi_master_awprot                                   (hps_0_h2f_lw_axi_master_awprot),                                          //                                                           .awprot
		.hps_0_h2f_lw_axi_master_awvalid                                  (hps_0_h2f_lw_axi_master_awvalid),                                         //                                                           .awvalid
		.hps_0_h2f_lw_axi_master_awready                                  (hps_0_h2f_lw_axi_master_awready),                                         //                                                           .awready
		.hps_0_h2f_lw_axi_master_wid                                      (hps_0_h2f_lw_axi_master_wid),                                             //                                                           .wid
		.hps_0_h2f_lw_axi_master_wdata                                    (hps_0_h2f_lw_axi_master_wdata),                                           //                                                           .wdata
		.hps_0_h2f_lw_axi_master_wstrb                                    (hps_0_h2f_lw_axi_master_wstrb),                                           //                                                           .wstrb
		.hps_0_h2f_lw_axi_master_wlast                                    (hps_0_h2f_lw_axi_master_wlast),                                           //                                                           .wlast
		.hps_0_h2f_lw_axi_master_wvalid                                   (hps_0_h2f_lw_axi_master_wvalid),                                          //                                                           .wvalid
		.hps_0_h2f_lw_axi_master_wready                                   (hps_0_h2f_lw_axi_master_wready),                                          //                                                           .wready
		.hps_0_h2f_lw_axi_master_bid                                      (hps_0_h2f_lw_axi_master_bid),                                             //                                                           .bid
		.hps_0_h2f_lw_axi_master_bresp                                    (hps_0_h2f_lw_axi_master_bresp),                                           //                                                           .bresp
		.hps_0_h2f_lw_axi_master_bvalid                                   (hps_0_h2f_lw_axi_master_bvalid),                                          //                                                           .bvalid
		.hps_0_h2f_lw_axi_master_bready                                   (hps_0_h2f_lw_axi_master_bready),                                          //                                                           .bready
		.hps_0_h2f_lw_axi_master_arid                                     (hps_0_h2f_lw_axi_master_arid),                                            //                                                           .arid
		.hps_0_h2f_lw_axi_master_araddr                                   (hps_0_h2f_lw_axi_master_araddr),                                          //                                                           .araddr
		.hps_0_h2f_lw_axi_master_arlen                                    (hps_0_h2f_lw_axi_master_arlen),                                           //                                                           .arlen
		.hps_0_h2f_lw_axi_master_arsize                                   (hps_0_h2f_lw_axi_master_arsize),                                          //                                                           .arsize
		.hps_0_h2f_lw_axi_master_arburst                                  (hps_0_h2f_lw_axi_master_arburst),                                         //                                                           .arburst
		.hps_0_h2f_lw_axi_master_arlock                                   (hps_0_h2f_lw_axi_master_arlock),                                          //                                                           .arlock
		.hps_0_h2f_lw_axi_master_arcache                                  (hps_0_h2f_lw_axi_master_arcache),                                         //                                                           .arcache
		.hps_0_h2f_lw_axi_master_arprot                                   (hps_0_h2f_lw_axi_master_arprot),                                          //                                                           .arprot
		.hps_0_h2f_lw_axi_master_arvalid                                  (hps_0_h2f_lw_axi_master_arvalid),                                         //                                                           .arvalid
		.hps_0_h2f_lw_axi_master_arready                                  (hps_0_h2f_lw_axi_master_arready),                                         //                                                           .arready
		.hps_0_h2f_lw_axi_master_rid                                      (hps_0_h2f_lw_axi_master_rid),                                             //                                                           .rid
		.hps_0_h2f_lw_axi_master_rdata                                    (hps_0_h2f_lw_axi_master_rdata),                                           //                                                           .rdata
		.hps_0_h2f_lw_axi_master_rresp                                    (hps_0_h2f_lw_axi_master_rresp),                                           //                                                           .rresp
		.hps_0_h2f_lw_axi_master_rlast                                    (hps_0_h2f_lw_axi_master_rlast),                                           //                                                           .rlast
		.hps_0_h2f_lw_axi_master_rvalid                                   (hps_0_h2f_lw_axi_master_rvalid),                                          //                                                           .rvalid
		.hps_0_h2f_lw_axi_master_rready                                   (hps_0_h2f_lw_axi_master_rready),                                          //                                                           .rready
		.clk_i_clk_clk                                                    (pll_0_sys_clk_clk),                                                       //                                                  clk_i_clk.clk
		.fpga_only_master_clk_reset_reset_bridge_in_reset_reset           (rst_controller_reset_out_reset),                                          //           fpga_only_master_clk_reset_reset_bridge_in_reset.reset
		.hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                                      // hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.nios2_qsys_0_reset_reset_bridge_in_reset_reset                   (rst_controller_reset_out_reset),                                          //                   nios2_qsys_0_reset_reset_bridge_in_reset.reset
		.sysid_reset_reset_bridge_in_reset_reset                          (rst_controller_001_reset_out_reset),                                      //                          sysid_reset_reset_bridge_in_reset.reset
		.fpga_only_master_master_address                                  (fpga_only_master_master_address),                                         //                                    fpga_only_master_master.address
		.fpga_only_master_master_waitrequest                              (fpga_only_master_master_waitrequest),                                     //                                                           .waitrequest
		.fpga_only_master_master_byteenable                               (fpga_only_master_master_byteenable),                                      //                                                           .byteenable
		.fpga_only_master_master_read                                     (fpga_only_master_master_read),                                            //                                                           .read
		.fpga_only_master_master_readdata                                 (fpga_only_master_master_readdata),                                        //                                                           .readdata
		.fpga_only_master_master_readdatavalid                            (fpga_only_master_master_readdatavalid),                                   //                                                           .readdatavalid
		.fpga_only_master_master_write                                    (fpga_only_master_master_write),                                           //                                                           .write
		.fpga_only_master_master_writedata                                (fpga_only_master_master_writedata),                                       //                                                           .writedata
		.nios2_qsys_0_data_master_address                                 (nios2_qsys_0_data_master_address),                                        //                                   nios2_qsys_0_data_master.address
		.nios2_qsys_0_data_master_waitrequest                             (nios2_qsys_0_data_master_waitrequest),                                    //                                                           .waitrequest
		.nios2_qsys_0_data_master_byteenable                              (nios2_qsys_0_data_master_byteenable),                                     //                                                           .byteenable
		.nios2_qsys_0_data_master_read                                    (nios2_qsys_0_data_master_read),                                           //                                                           .read
		.nios2_qsys_0_data_master_readdata                                (nios2_qsys_0_data_master_readdata),                                       //                                                           .readdata
		.nios2_qsys_0_data_master_write                                   (nios2_qsys_0_data_master_write),                                          //                                                           .write
		.nios2_qsys_0_data_master_writedata                               (nios2_qsys_0_data_master_writedata),                                      //                                                           .writedata
		.nios2_qsys_0_data_master_debugaccess                             (nios2_qsys_0_data_master_debugaccess),                                    //                                                           .debugaccess
		.nios2_qsys_0_instruction_master_address                          (nios2_qsys_0_instruction_master_address),                                 //                            nios2_qsys_0_instruction_master.address
		.nios2_qsys_0_instruction_master_waitrequest                      (nios2_qsys_0_instruction_master_waitrequest),                             //                                                           .waitrequest
		.nios2_qsys_0_instruction_master_read                             (nios2_qsys_0_instruction_master_read),                                    //                                                           .read
		.nios2_qsys_0_instruction_master_readdata                         (nios2_qsys_0_instruction_master_readdata),                                //                                                           .readdata
		.nios2_qsys_0_instruction_master_readdatavalid                    (nios2_qsys_0_instruction_master_readdatavalid),                           //                                                           .readdatavalid
		.avalon2fpga_slave_0_s1_address                                   (mm_interconnect_0_avalon2fpga_slave_0_s1_address),                        //                                     avalon2fpga_slave_0_s1.address
		.avalon2fpga_slave_0_s1_write                                     (mm_interconnect_0_avalon2fpga_slave_0_s1_write),                          //                                                           .write
		.avalon2fpga_slave_0_s1_read                                      (mm_interconnect_0_avalon2fpga_slave_0_s1_read),                           //                                                           .read
		.avalon2fpga_slave_0_s1_readdata                                  (mm_interconnect_0_avalon2fpga_slave_0_s1_readdata),                       //                                                           .readdata
		.avalon2fpga_slave_0_s1_writedata                                 (mm_interconnect_0_avalon2fpga_slave_0_s1_writedata),                      //                                                           .writedata
		.avalon2fpga_slave_0_s1_waitrequest                               (mm_interconnect_0_avalon2fpga_slave_0_s1_waitrequest),                    //                                                           .waitrequest
		.avalon_spi_amc7891_1_s1_address                                  (mm_interconnect_0_avalon_spi_amc7891_1_s1_address),                       //                                    avalon_spi_amc7891_1_s1.address
		.avalon_spi_amc7891_1_s1_write                                    (mm_interconnect_0_avalon_spi_amc7891_1_s1_write),                         //                                                           .write
		.avalon_spi_amc7891_1_s1_read                                     (mm_interconnect_0_avalon_spi_amc7891_1_s1_read),                          //                                                           .read
		.avalon_spi_amc7891_1_s1_readdata                                 (mm_interconnect_0_avalon_spi_amc7891_1_s1_readdata),                      //                                                           .readdata
		.avalon_spi_amc7891_1_s1_writedata                                (mm_interconnect_0_avalon_spi_amc7891_1_s1_writedata),                     //                                                           .writedata
		.avalon_spi_amc7891_1_s1_waitrequest                              (mm_interconnect_0_avalon_spi_amc7891_1_s1_waitrequest),                   //                                                           .waitrequest
		.avalon_spi_max31865_0_s1_address                                 (mm_interconnect_0_avalon_spi_max31865_0_s1_address),                      //                                   avalon_spi_max31865_0_s1.address
		.avalon_spi_max31865_0_s1_write                                   (mm_interconnect_0_avalon_spi_max31865_0_s1_write),                        //                                                           .write
		.avalon_spi_max31865_0_s1_read                                    (mm_interconnect_0_avalon_spi_max31865_0_s1_read),                         //                                                           .read
		.avalon_spi_max31865_0_s1_readdata                                (mm_interconnect_0_avalon_spi_max31865_0_s1_readdata),                     //                                                           .readdata
		.avalon_spi_max31865_0_s1_writedata                               (mm_interconnect_0_avalon_spi_max31865_0_s1_writedata),                    //                                                           .writedata
		.avalon_spi_max31865_0_s1_waitrequest                             (mm_interconnect_0_avalon_spi_max31865_0_s1_waitrequest),                  //                                                           .waitrequest
		.avalon_spi_max31865_1_s1_address                                 (mm_interconnect_0_avalon_spi_max31865_1_s1_address),                      //                                   avalon_spi_max31865_1_s1.address
		.avalon_spi_max31865_1_s1_write                                   (mm_interconnect_0_avalon_spi_max31865_1_s1_write),                        //                                                           .write
		.avalon_spi_max31865_1_s1_read                                    (mm_interconnect_0_avalon_spi_max31865_1_s1_read),                         //                                                           .read
		.avalon_spi_max31865_1_s1_readdata                                (mm_interconnect_0_avalon_spi_max31865_1_s1_readdata),                     //                                                           .readdata
		.avalon_spi_max31865_1_s1_writedata                               (mm_interconnect_0_avalon_spi_max31865_1_s1_writedata),                    //                                                           .writedata
		.avalon_spi_max31865_1_s1_waitrequest                             (mm_interconnect_0_avalon_spi_max31865_1_s1_waitrequest),                  //                                                           .waitrequest
		.avalon_spi_max31865_2_s1_address                                 (mm_interconnect_0_avalon_spi_max31865_2_s1_address),                      //                                   avalon_spi_max31865_2_s1.address
		.avalon_spi_max31865_2_s1_write                                   (mm_interconnect_0_avalon_spi_max31865_2_s1_write),                        //                                                           .write
		.avalon_spi_max31865_2_s1_read                                    (mm_interconnect_0_avalon_spi_max31865_2_s1_read),                         //                                                           .read
		.avalon_spi_max31865_2_s1_readdata                                (mm_interconnect_0_avalon_spi_max31865_2_s1_readdata),                     //                                                           .readdata
		.avalon_spi_max31865_2_s1_writedata                               (mm_interconnect_0_avalon_spi_max31865_2_s1_writedata),                    //                                                           .writedata
		.avalon_spi_max31865_2_s1_waitrequest                             (mm_interconnect_0_avalon_spi_max31865_2_s1_waitrequest),                  //                                                           .waitrequest
		.avalon_spi_max31865_3_s1_address                                 (mm_interconnect_0_avalon_spi_max31865_3_s1_address),                      //                                   avalon_spi_max31865_3_s1.address
		.avalon_spi_max31865_3_s1_write                                   (mm_interconnect_0_avalon_spi_max31865_3_s1_write),                        //                                                           .write
		.avalon_spi_max31865_3_s1_read                                    (mm_interconnect_0_avalon_spi_max31865_3_s1_read),                         //                                                           .read
		.avalon_spi_max31865_3_s1_readdata                                (mm_interconnect_0_avalon_spi_max31865_3_s1_readdata),                     //                                                           .readdata
		.avalon_spi_max31865_3_s1_writedata                               (mm_interconnect_0_avalon_spi_max31865_3_s1_writedata),                    //                                                           .writedata
		.avalon_spi_max31865_3_s1_waitrequest                             (mm_interconnect_0_avalon_spi_max31865_3_s1_waitrequest),                  //                                                           .waitrequest
		.avalon_spi_max31865_4_s1_address                                 (mm_interconnect_0_avalon_spi_max31865_4_s1_address),                      //                                   avalon_spi_max31865_4_s1.address
		.avalon_spi_max31865_4_s1_write                                   (mm_interconnect_0_avalon_spi_max31865_4_s1_write),                        //                                                           .write
		.avalon_spi_max31865_4_s1_read                                    (mm_interconnect_0_avalon_spi_max31865_4_s1_read),                         //                                                           .read
		.avalon_spi_max31865_4_s1_readdata                                (mm_interconnect_0_avalon_spi_max31865_4_s1_readdata),                     //                                                           .readdata
		.avalon_spi_max31865_4_s1_writedata                               (mm_interconnect_0_avalon_spi_max31865_4_s1_writedata),                    //                                                           .writedata
		.avalon_spi_max31865_4_s1_waitrequest                             (mm_interconnect_0_avalon_spi_max31865_4_s1_waitrequest),                  //                                                           .waitrequest
		.avalon_spi_max31865_5_s1_address                                 (mm_interconnect_0_avalon_spi_max31865_5_s1_address),                      //                                   avalon_spi_max31865_5_s1.address
		.avalon_spi_max31865_5_s1_write                                   (mm_interconnect_0_avalon_spi_max31865_5_s1_write),                        //                                                           .write
		.avalon_spi_max31865_5_s1_read                                    (mm_interconnect_0_avalon_spi_max31865_5_s1_read),                         //                                                           .read
		.avalon_spi_max31865_5_s1_readdata                                (mm_interconnect_0_avalon_spi_max31865_5_s1_readdata),                     //                                                           .readdata
		.avalon_spi_max31865_5_s1_writedata                               (mm_interconnect_0_avalon_spi_max31865_5_s1_writedata),                    //                                                           .writedata
		.avalon_spi_max31865_5_s1_waitrequest                             (mm_interconnect_0_avalon_spi_max31865_5_s1_waitrequest),                  //                                                           .waitrequest
		.flush_pump_pwm_duty_cycle_s1_address                             (mm_interconnect_0_flush_pump_pwm_duty_cycle_s1_address),                  //                               flush_pump_pwm_duty_cycle_s1.address
		.flush_pump_pwm_duty_cycle_s1_write                               (mm_interconnect_0_flush_pump_pwm_duty_cycle_s1_write),                    //                                                           .write
		.flush_pump_pwm_duty_cycle_s1_readdata                            (mm_interconnect_0_flush_pump_pwm_duty_cycle_s1_readdata),                 //                                                           .readdata
		.flush_pump_pwm_duty_cycle_s1_writedata                           (mm_interconnect_0_flush_pump_pwm_duty_cycle_s1_writedata),                //                                                           .writedata
		.flush_pump_pwm_duty_cycle_s1_chipselect                          (mm_interconnect_0_flush_pump_pwm_duty_cycle_s1_chipselect),               //                                                           .chipselect
		.flush_pump_pwm_freq_s1_address                                   (mm_interconnect_0_flush_pump_pwm_freq_s1_address),                        //                                     flush_pump_pwm_freq_s1.address
		.flush_pump_pwm_freq_s1_write                                     (mm_interconnect_0_flush_pump_pwm_freq_s1_write),                          //                                                           .write
		.flush_pump_pwm_freq_s1_readdata                                  (mm_interconnect_0_flush_pump_pwm_freq_s1_readdata),                       //                                                           .readdata
		.flush_pump_pwm_freq_s1_writedata                                 (mm_interconnect_0_flush_pump_pwm_freq_s1_writedata),                      //                                                           .writedata
		.flush_pump_pwm_freq_s1_chipselect                                (mm_interconnect_0_flush_pump_pwm_freq_s1_chipselect),                     //                                                           .chipselect
		.i2c_master_d_avalon_slave_address                                (mm_interconnect_0_i2c_master_d_avalon_slave_address),                     //                                  i2c_master_d_avalon_slave.address
		.i2c_master_d_avalon_slave_write                                  (mm_interconnect_0_i2c_master_d_avalon_slave_write),                       //                                                           .write
		.i2c_master_d_avalon_slave_readdata                               (mm_interconnect_0_i2c_master_d_avalon_slave_readdata),                    //                                                           .readdata
		.i2c_master_d_avalon_slave_writedata                              (mm_interconnect_0_i2c_master_d_avalon_slave_writedata),                   //                                                           .writedata
		.i2c_master_d_avalon_slave_waitrequest                            (~mm_interconnect_0_i2c_master_d_avalon_slave_waitrequest),                //                                                           .waitrequest
		.i2c_master_d_avalon_slave_chipselect                             (mm_interconnect_0_i2c_master_d_avalon_slave_chipselect),                  //                                                           .chipselect
		.i2c_master_f_avalon_slave_address                                (mm_interconnect_0_i2c_master_f_avalon_slave_address),                     //                                  i2c_master_f_avalon_slave.address
		.i2c_master_f_avalon_slave_write                                  (mm_interconnect_0_i2c_master_f_avalon_slave_write),                       //                                                           .write
		.i2c_master_f_avalon_slave_readdata                               (mm_interconnect_0_i2c_master_f_avalon_slave_readdata),                    //                                                           .readdata
		.i2c_master_f_avalon_slave_writedata                              (mm_interconnect_0_i2c_master_f_avalon_slave_writedata),                   //                                                           .writedata
		.i2c_master_f_avalon_slave_waitrequest                            (~mm_interconnect_0_i2c_master_f_avalon_slave_waitrequest),                //                                                           .waitrequest
		.i2c_master_f_avalon_slave_chipselect                             (mm_interconnect_0_i2c_master_f_avalon_slave_chipselect),                  //                                                           .chipselect
		.i2c_master_is1_avalon_slave_address                              (mm_interconnect_0_i2c_master_is1_avalon_slave_address),                   //                                i2c_master_is1_avalon_slave.address
		.i2c_master_is1_avalon_slave_write                                (mm_interconnect_0_i2c_master_is1_avalon_slave_write),                     //                                                           .write
		.i2c_master_is1_avalon_slave_readdata                             (mm_interconnect_0_i2c_master_is1_avalon_slave_readdata),                  //                                                           .readdata
		.i2c_master_is1_avalon_slave_writedata                            (mm_interconnect_0_i2c_master_is1_avalon_slave_writedata),                 //                                                           .writedata
		.i2c_master_is1_avalon_slave_waitrequest                          (~mm_interconnect_0_i2c_master_is1_avalon_slave_waitrequest),              //                                                           .waitrequest
		.i2c_master_is1_avalon_slave_chipselect                           (mm_interconnect_0_i2c_master_is1_avalon_slave_chipselect),                //                                                           .chipselect
		.i2c_master_is2_avalon_slave_address                              (mm_interconnect_0_i2c_master_is2_avalon_slave_address),                   //                                i2c_master_is2_avalon_slave.address
		.i2c_master_is2_avalon_slave_write                                (mm_interconnect_0_i2c_master_is2_avalon_slave_write),                     //                                                           .write
		.i2c_master_is2_avalon_slave_readdata                             (mm_interconnect_0_i2c_master_is2_avalon_slave_readdata),                  //                                                           .readdata
		.i2c_master_is2_avalon_slave_writedata                            (mm_interconnect_0_i2c_master_is2_avalon_slave_writedata),                 //                                                           .writedata
		.i2c_master_is2_avalon_slave_waitrequest                          (~mm_interconnect_0_i2c_master_is2_avalon_slave_waitrequest),              //                                                           .waitrequest
		.i2c_master_is2_avalon_slave_chipselect                           (mm_interconnect_0_i2c_master_is2_avalon_slave_chipselect),                //                                                           .chipselect
		.i2c_master_is3_avalon_slave_address                              (mm_interconnect_0_i2c_master_is3_avalon_slave_address),                   //                                i2c_master_is3_avalon_slave.address
		.i2c_master_is3_avalon_slave_write                                (mm_interconnect_0_i2c_master_is3_avalon_slave_write),                     //                                                           .write
		.i2c_master_is3_avalon_slave_readdata                             (mm_interconnect_0_i2c_master_is3_avalon_slave_readdata),                  //                                                           .readdata
		.i2c_master_is3_avalon_slave_writedata                            (mm_interconnect_0_i2c_master_is3_avalon_slave_writedata),                 //                                                           .writedata
		.i2c_master_is3_avalon_slave_waitrequest                          (~mm_interconnect_0_i2c_master_is3_avalon_slave_waitrequest),              //                                                           .waitrequest
		.i2c_master_is3_avalon_slave_chipselect                           (mm_interconnect_0_i2c_master_is3_avalon_slave_chipselect),                //                                                           .chipselect
		.i2c_master_is4_avalon_slave_address                              (mm_interconnect_0_i2c_master_is4_avalon_slave_address),                   //                                i2c_master_is4_avalon_slave.address
		.i2c_master_is4_avalon_slave_write                                (mm_interconnect_0_i2c_master_is4_avalon_slave_write),                     //                                                           .write
		.i2c_master_is4_avalon_slave_readdata                             (mm_interconnect_0_i2c_master_is4_avalon_slave_readdata),                  //                                                           .readdata
		.i2c_master_is4_avalon_slave_writedata                            (mm_interconnect_0_i2c_master_is4_avalon_slave_writedata),                 //                                                           .writedata
		.i2c_master_is4_avalon_slave_waitrequest                          (~mm_interconnect_0_i2c_master_is4_avalon_slave_waitrequest),              //                                                           .waitrequest
		.i2c_master_is4_avalon_slave_chipselect                           (mm_interconnect_0_i2c_master_is4_avalon_slave_chipselect),                //                                                           .chipselect
		.i2c_master_p_avalon_slave_address                                (mm_interconnect_0_i2c_master_p_avalon_slave_address),                     //                                  i2c_master_p_avalon_slave.address
		.i2c_master_p_avalon_slave_write                                  (mm_interconnect_0_i2c_master_p_avalon_slave_write),                       //                                                           .write
		.i2c_master_p_avalon_slave_readdata                               (mm_interconnect_0_i2c_master_p_avalon_slave_readdata),                    //                                                           .readdata
		.i2c_master_p_avalon_slave_writedata                              (mm_interconnect_0_i2c_master_p_avalon_slave_writedata),                   //                                                           .writedata
		.i2c_master_p_avalon_slave_waitrequest                            (~mm_interconnect_0_i2c_master_p_avalon_slave_waitrequest),                //                                                           .waitrequest
		.i2c_master_p_avalon_slave_chipselect                             (mm_interconnect_0_i2c_master_p_avalon_slave_chipselect),                  //                                                           .chipselect
		.jtag_uart_avalon_jtag_slave_address                              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),                   //                                jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),                     //                                                           .write
		.jtag_uart_avalon_jtag_slave_read                                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),                      //                                                           .read
		.jtag_uart_avalon_jtag_slave_readdata                             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),                  //                                                           .readdata
		.jtag_uart_avalon_jtag_slave_writedata                            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),                 //                                                           .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),               //                                                           .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),                //                                                           .chipselect
		.nios2_qsys_0_debug_mem_slave_address                             (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_address),                  //                               nios2_qsys_0_debug_mem_slave.address
		.nios2_qsys_0_debug_mem_slave_write                               (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_write),                    //                                                           .write
		.nios2_qsys_0_debug_mem_slave_read                                (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_read),                     //                                                           .read
		.nios2_qsys_0_debug_mem_slave_readdata                            (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_readdata),                 //                                                           .readdata
		.nios2_qsys_0_debug_mem_slave_writedata                           (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_writedata),                //                                                           .writedata
		.nios2_qsys_0_debug_mem_slave_byteenable                          (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_byteenable),               //                                                           .byteenable
		.nios2_qsys_0_debug_mem_slave_waitrequest                         (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_waitrequest),              //                                                           .waitrequest
		.nios2_qsys_0_debug_mem_slave_debugaccess                         (mm_interconnect_0_nios2_qsys_0_debug_mem_slave_debugaccess),              //                                                           .debugaccess
		.onchip_memory_nios_arm_s1_address                                (mm_interconnect_0_onchip_memory_nios_arm_s1_address),                     //                                  onchip_memory_nios_arm_s1.address
		.onchip_memory_nios_arm_s1_write                                  (mm_interconnect_0_onchip_memory_nios_arm_s1_write),                       //                                                           .write
		.onchip_memory_nios_arm_s1_readdata                               (mm_interconnect_0_onchip_memory_nios_arm_s1_readdata),                    //                                                           .readdata
		.onchip_memory_nios_arm_s1_writedata                              (mm_interconnect_0_onchip_memory_nios_arm_s1_writedata),                   //                                                           .writedata
		.onchip_memory_nios_arm_s1_byteenable                             (mm_interconnect_0_onchip_memory_nios_arm_s1_byteenable),                  //                                                           .byteenable
		.onchip_memory_nios_arm_s1_chipselect                             (mm_interconnect_0_onchip_memory_nios_arm_s1_chipselect),                  //                                                           .chipselect
		.onchip_memory_nios_arm_s1_clken                                  (mm_interconnect_0_onchip_memory_nios_arm_s1_clken),                       //                                                           .clken
		.onchip_memory_nios_arm_s2_address                                (mm_interconnect_0_onchip_memory_nios_arm_s2_address),                     //                                  onchip_memory_nios_arm_s2.address
		.onchip_memory_nios_arm_s2_write                                  (mm_interconnect_0_onchip_memory_nios_arm_s2_write),                       //                                                           .write
		.onchip_memory_nios_arm_s2_readdata                               (mm_interconnect_0_onchip_memory_nios_arm_s2_readdata),                    //                                                           .readdata
		.onchip_memory_nios_arm_s2_writedata                              (mm_interconnect_0_onchip_memory_nios_arm_s2_writedata),                   //                                                           .writedata
		.onchip_memory_nios_arm_s2_byteenable                             (mm_interconnect_0_onchip_memory_nios_arm_s2_byteenable),                  //                                                           .byteenable
		.onchip_memory_nios_arm_s2_chipselect                             (mm_interconnect_0_onchip_memory_nios_arm_s2_chipselect),                  //                                                           .chipselect
		.onchip_memory_nios_arm_s2_clken                                  (mm_interconnect_0_onchip_memory_nios_arm_s2_clken),                       //                                                           .clken
		.onchip_memory_nios_cpu_s1_address                                (mm_interconnect_0_onchip_memory_nios_cpu_s1_address),                     //                                  onchip_memory_nios_cpu_s1.address
		.onchip_memory_nios_cpu_s1_write                                  (mm_interconnect_0_onchip_memory_nios_cpu_s1_write),                       //                                                           .write
		.onchip_memory_nios_cpu_s1_readdata                               (mm_interconnect_0_onchip_memory_nios_cpu_s1_readdata),                    //                                                           .readdata
		.onchip_memory_nios_cpu_s1_writedata                              (mm_interconnect_0_onchip_memory_nios_cpu_s1_writedata),                   //                                                           .writedata
		.onchip_memory_nios_cpu_s1_byteenable                             (mm_interconnect_0_onchip_memory_nios_cpu_s1_byteenable),                  //                                                           .byteenable
		.onchip_memory_nios_cpu_s1_chipselect                             (mm_interconnect_0_onchip_memory_nios_cpu_s1_chipselect),                  //                                                           .chipselect
		.onchip_memory_nios_cpu_s1_clken                                  (mm_interconnect_0_onchip_memory_nios_cpu_s1_clken),                       //                                                           .clken
		.onchip_memory_nios_cpu_s2_address                                (mm_interconnect_0_onchip_memory_nios_cpu_s2_address),                     //                                  onchip_memory_nios_cpu_s2.address
		.onchip_memory_nios_cpu_s2_write                                  (mm_interconnect_0_onchip_memory_nios_cpu_s2_write),                       //                                                           .write
		.onchip_memory_nios_cpu_s2_readdata                               (mm_interconnect_0_onchip_memory_nios_cpu_s2_readdata),                    //                                                           .readdata
		.onchip_memory_nios_cpu_s2_writedata                              (mm_interconnect_0_onchip_memory_nios_cpu_s2_writedata),                   //                                                           .writedata
		.onchip_memory_nios_cpu_s2_byteenable                             (mm_interconnect_0_onchip_memory_nios_cpu_s2_byteenable),                  //                                                           .byteenable
		.onchip_memory_nios_cpu_s2_chipselect                             (mm_interconnect_0_onchip_memory_nios_cpu_s2_chipselect),                  //                                                           .chipselect
		.onchip_memory_nios_cpu_s2_clken                                  (mm_interconnect_0_onchip_memory_nios_cpu_s2_clken),                       //                                                           .clken
		.pio_input_s1_address                                             (mm_interconnect_0_pio_input_s1_address),                                  //                                               pio_input_s1.address
		.pio_input_s1_write                                               (mm_interconnect_0_pio_input_s1_write),                                    //                                                           .write
		.pio_input_s1_readdata                                            (mm_interconnect_0_pio_input_s1_readdata),                                 //                                                           .readdata
		.pio_input_s1_writedata                                           (mm_interconnect_0_pio_input_s1_writedata),                                //                                                           .writedata
		.pio_input_s1_chipselect                                          (mm_interconnect_0_pio_input_s1_chipselect),                               //                                                           .chipselect
		.pio_output_s1_address                                            (mm_interconnect_0_pio_output_s1_address),                                 //                                              pio_output_s1.address
		.pio_output_s1_write                                              (mm_interconnect_0_pio_output_s1_write),                                   //                                                           .write
		.pio_output_s1_readdata                                           (mm_interconnect_0_pio_output_s1_readdata),                                //                                                           .readdata
		.pio_output_s1_writedata                                          (mm_interconnect_0_pio_output_s1_writedata),                               //                                                           .writedata
		.pio_output_s1_chipselect                                         (mm_interconnect_0_pio_output_s1_chipselect),                              //                                                           .chipselect
		.pio_reset_nios_s1_address                                        (mm_interconnect_0_pio_reset_nios_s1_address),                             //                                          pio_reset_nios_s1.address
		.pio_reset_nios_s1_write                                          (mm_interconnect_0_pio_reset_nios_s1_write),                               //                                                           .write
		.pio_reset_nios_s1_readdata                                       (mm_interconnect_0_pio_reset_nios_s1_readdata),                            //                                                           .readdata
		.pio_reset_nios_s1_writedata                                      (mm_interconnect_0_pio_reset_nios_s1_writedata),                           //                                                           .writedata
		.pio_reset_nios_s1_chipselect                                     (mm_interconnect_0_pio_reset_nios_s1_chipselect),                          //                                                           .chipselect
		.pio_watchdog_cnt_s1_address                                      (mm_interconnect_0_pio_watchdog_cnt_s1_address),                           //                                        pio_watchdog_cnt_s1.address
		.pio_watchdog_cnt_s1_write                                        (mm_interconnect_0_pio_watchdog_cnt_s1_write),                             //                                                           .write
		.pio_watchdog_cnt_s1_readdata                                     (mm_interconnect_0_pio_watchdog_cnt_s1_readdata),                          //                                                           .readdata
		.pio_watchdog_cnt_s1_writedata                                    (mm_interconnect_0_pio_watchdog_cnt_s1_writedata),                         //                                                           .writedata
		.pio_watchdog_cnt_s1_chipselect                                   (mm_interconnect_0_pio_watchdog_cnt_s1_chipselect),                        //                                                           .chipselect
		.pio_watchdog_freq_s1_address                                     (mm_interconnect_0_pio_watchdog_freq_s1_address),                          //                                       pio_watchdog_freq_s1.address
		.pio_watchdog_freq_s1_write                                       (mm_interconnect_0_pio_watchdog_freq_s1_write),                            //                                                           .write
		.pio_watchdog_freq_s1_readdata                                    (mm_interconnect_0_pio_watchdog_freq_s1_readdata),                         //                                                           .readdata
		.pio_watchdog_freq_s1_writedata                                   (mm_interconnect_0_pio_watchdog_freq_s1_writedata),                        //                                                           .writedata
		.pio_watchdog_freq_s1_chipselect                                  (mm_interconnect_0_pio_watchdog_freq_s1_chipselect),                       //                                                           .chipselect
		.sysid_control_slave_address                                      (mm_interconnect_0_sysid_control_slave_address),                           //                                        sysid_control_slave.address
		.sysid_control_slave_readdata                                     (mm_interconnect_0_sysid_control_slave_readdata),                          //                                                           .readdata
		.timer_0_s1_address                                               (mm_interconnect_0_timer_0_s1_address),                                    //                                                 timer_0_s1.address
		.timer_0_s1_write                                                 (mm_interconnect_0_timer_0_s1_write),                                      //                                                           .write
		.timer_0_s1_readdata                                              (mm_interconnect_0_timer_0_s1_readdata),                                   //                                                           .readdata
		.timer_0_s1_writedata                                             (mm_interconnect_0_timer_0_s1_writedata),                                  //                                                           .writedata
		.timer_0_s1_chipselect                                            (mm_interconnect_0_timer_0_s1_chipselect),                                 //                                                           .chipselect
		.timer_1_s1_address                                               (mm_interconnect_0_timer_1_s1_address),                                    //                                                 timer_1_s1.address
		.timer_1_s1_write                                                 (mm_interconnect_0_timer_1_s1_write),                                      //                                                           .write
		.timer_1_s1_readdata                                              (mm_interconnect_0_timer_1_s1_readdata),                                   //                                                           .readdata
		.timer_1_s1_writedata                                             (mm_interconnect_0_timer_1_s1_writedata),                                  //                                                           .writedata
		.timer_1_s1_chipselect                                            (mm_interconnect_0_timer_1_s1_chipselect),                                 //                                                           .chipselect
		.timer_2_s1_address                                               (mm_interconnect_0_timer_2_s1_address),                                    //                                                 timer_2_s1.address
		.timer_2_s1_write                                                 (mm_interconnect_0_timer_2_s1_write),                                      //                                                           .write
		.timer_2_s1_readdata                                              (mm_interconnect_0_timer_2_s1_readdata),                                   //                                                           .readdata
		.timer_2_s1_writedata                                             (mm_interconnect_0_timer_2_s1_writedata),                                  //                                                           .writedata
		.timer_2_s1_chipselect                                            (mm_interconnect_0_timer_2_s1_chipselect)                                  //                                                           .chipselect
	);

	fluid_board_soc_irq_mapper irq_mapper (
		.clk           (),                         //       clk.clk
		.reset         (),                         // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq), // receiver0.irq
		.sender_irq    (hps_0_f2h_irq0_irq)        //    sender.irq
	);

	fluid_board_soc_irq_mapper_001 irq_mapper_001 (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq1_irq)  //    sender.irq
	);

	fluid_board_soc_irq_mapper_002 irq_mapper_002 (
		.clk            (pll_0_sys_clk_clk),              //        clk.clk
		.reset          (rst_controller_reset_out_reset), //  clk_reset.reset
		.receiver0_irq  (irq_mapper_002_receiver0_irq),   //  receiver0.irq
		.receiver1_irq  (irq_mapper_002_receiver1_irq),   //  receiver1.irq
		.receiver2_irq  (irq_mapper_002_receiver2_irq),   //  receiver2.irq
		.receiver3_irq  (irq_mapper_002_receiver3_irq),   //  receiver3.irq
		.receiver4_irq  (irq_mapper_002_receiver4_irq),   //  receiver4.irq
		.receiver5_irq  (irq_mapper_002_receiver5_irq),   //  receiver5.irq
		.receiver6_irq  (irq_mapper_002_receiver6_irq),   //  receiver6.irq
		.receiver7_irq  (irq_mapper_002_receiver7_irq),   //  receiver7.irq
		.receiver8_irq  (irq_mapper_002_receiver8_irq),   //  receiver8.irq
		.receiver9_irq  (irq_mapper_002_receiver9_irq),   //  receiver9.irq
		.receiver10_irq (irq_mapper_receiver0_irq),       // receiver10.irq
		.receiver11_irq (irq_mapper_002_receiver11_irq),  // receiver11.irq
		.sender_irq     (nios2_qsys_0_irq_irq)            //     sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~qsys_reset_reset_n),                // reset_in0.reset
		.clk            (pll_0_sys_clk_clk),                  //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~qsys_reset_reset_n),                    // reset_in0.reset
		.reset_in1      (~hps_0_h2f_reset_reset),                 // reset_in1.reset
		.clk            (pll_0_sys_clk_clk),                      //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.clk            (pll_0_sys_clk_clk),                  //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	assign pll_0_sys_reset_reset_n = qsys_reset_reset_n;

endmodule
