-- fluid_board_soc.vhd

-- Generated using ACDS version 14.0 200 at 2015.12.23.13:39:17

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity fluid_board_soc is
	port (
		hps_io_hps_io_emac0_inst_TX_CLK                    : out   std_logic;                                        --                                hps_io.hps_io_emac0_inst_TX_CLK
		hps_io_hps_io_emac0_inst_TXD0                      : out   std_logic;                                        --                                      .hps_io_emac0_inst_TXD0
		hps_io_hps_io_emac0_inst_TXD1                      : out   std_logic;                                        --                                      .hps_io_emac0_inst_TXD1
		hps_io_hps_io_emac0_inst_TXD2                      : out   std_logic;                                        --                                      .hps_io_emac0_inst_TXD2
		hps_io_hps_io_emac0_inst_TXD3                      : out   std_logic;                                        --                                      .hps_io_emac0_inst_TXD3
		hps_io_hps_io_emac0_inst_RXD0                      : in    std_logic                     := '0';             --                                      .hps_io_emac0_inst_RXD0
		hps_io_hps_io_emac0_inst_MDIO                      : inout std_logic                     := '0';             --                                      .hps_io_emac0_inst_MDIO
		hps_io_hps_io_emac0_inst_MDC                       : out   std_logic;                                        --                                      .hps_io_emac0_inst_MDC
		hps_io_hps_io_emac0_inst_RX_CTL                    : in    std_logic                     := '0';             --                                      .hps_io_emac0_inst_RX_CTL
		hps_io_hps_io_emac0_inst_TX_CTL                    : out   std_logic;                                        --                                      .hps_io_emac0_inst_TX_CTL
		hps_io_hps_io_emac0_inst_RX_CLK                    : in    std_logic                     := '0';             --                                      .hps_io_emac0_inst_RX_CLK
		hps_io_hps_io_emac0_inst_RXD1                      : in    std_logic                     := '0';             --                                      .hps_io_emac0_inst_RXD1
		hps_io_hps_io_emac0_inst_RXD2                      : in    std_logic                     := '0';             --                                      .hps_io_emac0_inst_RXD2
		hps_io_hps_io_emac0_inst_RXD3                      : in    std_logic                     := '0';             --                                      .hps_io_emac0_inst_RXD3
		hps_io_hps_io_uart0_inst_RX                        : in    std_logic                     := '0';             --                                      .hps_io_uart0_inst_RX
		hps_io_hps_io_uart0_inst_TX                        : out   std_logic;                                        --                                      .hps_io_uart0_inst_TX
		hps_io_hps_io_gpio_inst_GPIO26                     : inout std_logic                     := '0';             --                                      .hps_io_gpio_inst_GPIO26
		hps_io_hps_io_gpio_inst_GPIO28                     : inout std_logic                     := '0';             --                                      .hps_io_gpio_inst_GPIO28
		hps_io_hps_io_gpio_inst_GPIO59                     : inout std_logic                     := '0';             --                                      .hps_io_gpio_inst_GPIO59
		memory_mem_a                                       : out   std_logic_vector(14 downto 0);                    --                                memory.mem_a
		memory_mem_ba                                      : out   std_logic_vector(2 downto 0);                     --                                      .mem_ba
		memory_mem_ck                                      : out   std_logic;                                        --                                      .mem_ck
		memory_mem_ck_n                                    : out   std_logic;                                        --                                      .mem_ck_n
		memory_mem_cke                                     : out   std_logic;                                        --                                      .mem_cke
		memory_mem_cs_n                                    : out   std_logic;                                        --                                      .mem_cs_n
		memory_mem_ras_n                                   : out   std_logic;                                        --                                      .mem_ras_n
		memory_mem_cas_n                                   : out   std_logic;                                        --                                      .mem_cas_n
		memory_mem_we_n                                    : out   std_logic;                                        --                                      .mem_we_n
		memory_mem_reset_n                                 : out   std_logic;                                        --                                      .mem_reset_n
		memory_mem_dq                                      : inout std_logic_vector(31 downto 0) := (others => '0'); --                                      .mem_dq
		memory_mem_dqs                                     : inout std_logic_vector(3 downto 0)  := (others => '0'); --                                      .mem_dqs
		memory_mem_dqs_n                                   : inout std_logic_vector(3 downto 0)  := (others => '0'); --                                      .mem_dqs_n
		memory_mem_odt                                     : out   std_logic;                                        --                                      .mem_odt
		memory_mem_dm                                      : out   std_logic_vector(3 downto 0);                     --                                      .mem_dm
		memory_oct_rzqin                                   : in    std_logic                     := '0';             --                                      .oct_rzqin
		hps_0_uart1_cts                                    : in    std_logic                     := '0';             --                           hps_0_uart1.cts
		hps_0_uart1_dsr                                    : in    std_logic                     := '0';             --                                      .dsr
		hps_0_uart1_dcd                                    : in    std_logic                     := '0';             --                                      .dcd
		hps_0_uart1_ri                                     : in    std_logic                     := '0';             --                                      .ri
		hps_0_uart1_dtr                                    : out   std_logic;                                        --                                      .dtr
		hps_0_uart1_rts                                    : out   std_logic;                                        --                                      .rts
		hps_0_uart1_out1_n                                 : out   std_logic;                                        --                                      .out1_n
		hps_0_uart1_out2_n                                 : out   std_logic;                                        --                                      .out2_n
		hps_0_uart1_rxd                                    : in    std_logic                     := '0';             --                                      .rxd
		hps_0_uart1_txd                                    : out   std_logic;                                        --                                      .txd
		pll_0_locked_export                                : out   std_logic;                                        --                          pll_0_locked.export
		pll_0_reset_reset                                  : in    std_logic                     := '0';             --                           pll_0_reset.reset
		pll_0_sys_clk_clk                                  : out   std_logic;                                        --                         pll_0_sys_clk.clk
		pll_0_refclk_clk                                   : in    std_logic                     := '0';             --                          pll_0_refclk.clk
		qsys_reset_reset_n                                 : in    std_logic                     := '0';             --                            qsys_reset.reset_n
		pll_0_sys_reset_reset_n                            : out   std_logic;                                        --                       pll_0_sys_reset.reset_n
		i2c_master_is4_conduit_end_scl                     : inout std_logic                     := '0';             --            i2c_master_is4_conduit_end.scl
		i2c_master_is4_conduit_end_sda                     : inout std_logic                     := '0';             --                                      .sda
		i2c_master_is1_conduit_end_scl                     : inout std_logic                     := '0';             --            i2c_master_is1_conduit_end.scl
		i2c_master_is1_conduit_end_sda                     : inout std_logic                     := '0';             --                                      .sda
		i2c_master_is2_conduit_end_scl                     : inout std_logic                     := '0';             --            i2c_master_is2_conduit_end.scl
		i2c_master_is2_conduit_end_sda                     : inout std_logic                     := '0';             --                                      .sda
		i2c_master_is3_conduit_end_scl                     : inout std_logic                     := '0';             --            i2c_master_is3_conduit_end.scl
		i2c_master_is3_conduit_end_sda                     : inout std_logic                     := '0';             --                                      .sda
		nios2_qsys_0_cpu_resetrequest_conduit_resetrequest : in    std_logic                     := '0';             -- nios2_qsys_0_cpu_resetrequest_conduit.resetrequest
		nios2_qsys_0_cpu_resetrequest_conduit_resettaken   : out   std_logic;                                        --                                      .resettaken
		pio_input_external_connection_export               : in    std_logic_vector(3 downto 0)  := (others => '0'); --         pio_input_external_connection.export
		pio_output_external_connection_export              : out   std_logic_vector(7 downto 0);                     --        pio_output_external_connection.export
		i2c_master_d_conduit_end_scl                       : inout std_logic                     := '0';             --              i2c_master_d_conduit_end.scl
		i2c_master_d_conduit_end_sda                       : inout std_logic                     := '0';             --                                      .sda
		i2c_master_f_conduit_end_scl                       : inout std_logic                     := '0';             --              i2c_master_f_conduit_end.scl
		i2c_master_f_conduit_end_sda                       : inout std_logic                     := '0';             --                                      .sda
		i2c_master_p_conduit_end_scl                       : inout std_logic                     := '0';             --              i2c_master_p_conduit_end.scl
		i2c_master_p_conduit_end_sda                       : inout std_logic                     := '0';             --                                      .sda
		pio_reset_nios_external_connection_export          : out   std_logic;                                        --    pio_reset_nios_external_connection.export
		avalon_spi_amc7891_1_conduit_end_sclk              : out   std_logic;                                        --      avalon_spi_amc7891_1_conduit_end.sclk
		avalon_spi_amc7891_1_conduit_end_cs_n              : out   std_logic;                                        --                                      .cs_n
		avalon_spi_amc7891_1_conduit_end_sdio              : out   std_logic;                                        --                                      .sdio
		avalon_spi_amc7891_1_conduit_end_sdo               : in    std_logic                     := '0';             --                                      .sdo
		avalon_spi_amc7891_0_conduit_end_sclk              : out   std_logic;                                        --      avalon_spi_amc7891_0_conduit_end.sclk
		avalon_spi_amc7891_0_conduit_end_cs_n              : out   std_logic;                                        --                                      .cs_n
		avalon_spi_amc7891_0_conduit_end_sdio              : out   std_logic;                                        --                                      .sdio
		avalon_spi_amc7891_0_conduit_end_sdo               : in    std_logic                     := '0'              --                                      .sdo
	);
end entity fluid_board_soc;

architecture rtl of fluid_board_soc is
	component fluid_board_soc_hps_0 is
		generic (
			F2S_Width : integer := 2;
			S2F_Width : integer := 2
		);
		port (
			uart1_cts                : in    std_logic                     := 'X';             -- cts
			uart1_dsr                : in    std_logic                     := 'X';             -- dsr
			uart1_dcd                : in    std_logic                     := 'X';             -- dcd
			uart1_ri                 : in    std_logic                     := 'X';             -- ri
			uart1_dtr                : out   std_logic;                                        -- dtr
			uart1_rts                : out   std_logic;                                        -- rts
			uart1_out1_n             : out   std_logic;                                        -- out1_n
			uart1_out2_n             : out   std_logic;                                        -- out2_n
			uart1_rxd                : in    std_logic                     := 'X';             -- rxd
			uart1_txd                : out   std_logic;                                        -- txd
			mem_a                    : out   std_logic_vector(14 downto 0);                    -- mem_a
			mem_ba                   : out   std_logic_vector(2 downto 0);                     -- mem_ba
			mem_ck                   : out   std_logic;                                        -- mem_ck
			mem_ck_n                 : out   std_logic;                                        -- mem_ck_n
			mem_cke                  : out   std_logic;                                        -- mem_cke
			mem_cs_n                 : out   std_logic;                                        -- mem_cs_n
			mem_ras_n                : out   std_logic;                                        -- mem_ras_n
			mem_cas_n                : out   std_logic;                                        -- mem_cas_n
			mem_we_n                 : out   std_logic;                                        -- mem_we_n
			mem_reset_n              : out   std_logic;                                        -- mem_reset_n
			mem_dq                   : inout std_logic_vector(31 downto 0) := (others => 'X'); -- mem_dq
			mem_dqs                  : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs
			mem_dqs_n                : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs_n
			mem_odt                  : out   std_logic;                                        -- mem_odt
			mem_dm                   : out   std_logic_vector(3 downto 0);                     -- mem_dm
			oct_rzqin                : in    std_logic                     := 'X';             -- oct_rzqin
			hps_io_emac0_inst_TX_CLK : out   std_logic;                                        -- hps_io_emac0_inst_TX_CLK
			hps_io_emac0_inst_TXD0   : out   std_logic;                                        -- hps_io_emac0_inst_TXD0
			hps_io_emac0_inst_TXD1   : out   std_logic;                                        -- hps_io_emac0_inst_TXD1
			hps_io_emac0_inst_TXD2   : out   std_logic;                                        -- hps_io_emac0_inst_TXD2
			hps_io_emac0_inst_TXD3   : out   std_logic;                                        -- hps_io_emac0_inst_TXD3
			hps_io_emac0_inst_RXD0   : in    std_logic                     := 'X';             -- hps_io_emac0_inst_RXD0
			hps_io_emac0_inst_MDIO   : inout std_logic                     := 'X';             -- hps_io_emac0_inst_MDIO
			hps_io_emac0_inst_MDC    : out   std_logic;                                        -- hps_io_emac0_inst_MDC
			hps_io_emac0_inst_RX_CTL : in    std_logic                     := 'X';             -- hps_io_emac0_inst_RX_CTL
			hps_io_emac0_inst_TX_CTL : out   std_logic;                                        -- hps_io_emac0_inst_TX_CTL
			hps_io_emac0_inst_RX_CLK : in    std_logic                     := 'X';             -- hps_io_emac0_inst_RX_CLK
			hps_io_emac0_inst_RXD1   : in    std_logic                     := 'X';             -- hps_io_emac0_inst_RXD1
			hps_io_emac0_inst_RXD2   : in    std_logic                     := 'X';             -- hps_io_emac0_inst_RXD2
			hps_io_emac0_inst_RXD3   : in    std_logic                     := 'X';             -- hps_io_emac0_inst_RXD3
			hps_io_uart0_inst_RX     : in    std_logic                     := 'X';             -- hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX     : out   std_logic;                                        -- hps_io_uart0_inst_TX
			hps_io_gpio_inst_GPIO26  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO26
			hps_io_gpio_inst_GPIO28  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO28
			hps_io_gpio_inst_GPIO59  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO59
			h2f_rst_n                : out   std_logic;                                        -- reset_n
			h2f_axi_clk              : in    std_logic                     := 'X';             -- clk
			h2f_AWID                 : out   std_logic_vector(11 downto 0);                    -- awid
			h2f_AWADDR               : out   std_logic_vector(29 downto 0);                    -- awaddr
			h2f_AWLEN                : out   std_logic_vector(3 downto 0);                     -- awlen
			h2f_AWSIZE               : out   std_logic_vector(2 downto 0);                     -- awsize
			h2f_AWBURST              : out   std_logic_vector(1 downto 0);                     -- awburst
			h2f_AWLOCK               : out   std_logic_vector(1 downto 0);                     -- awlock
			h2f_AWCACHE              : out   std_logic_vector(3 downto 0);                     -- awcache
			h2f_AWPROT               : out   std_logic_vector(2 downto 0);                     -- awprot
			h2f_AWVALID              : out   std_logic;                                        -- awvalid
			h2f_AWREADY              : in    std_logic                     := 'X';             -- awready
			h2f_WID                  : out   std_logic_vector(11 downto 0);                    -- wid
			h2f_WDATA                : out   std_logic_vector(63 downto 0);                    -- wdata
			h2f_WSTRB                : out   std_logic_vector(7 downto 0);                     -- wstrb
			h2f_WLAST                : out   std_logic;                                        -- wlast
			h2f_WVALID               : out   std_logic;                                        -- wvalid
			h2f_WREADY               : in    std_logic                     := 'X';             -- wready
			h2f_BID                  : in    std_logic_vector(11 downto 0) := (others => 'X'); -- bid
			h2f_BRESP                : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			h2f_BVALID               : in    std_logic                     := 'X';             -- bvalid
			h2f_BREADY               : out   std_logic;                                        -- bready
			h2f_ARID                 : out   std_logic_vector(11 downto 0);                    -- arid
			h2f_ARADDR               : out   std_logic_vector(29 downto 0);                    -- araddr
			h2f_ARLEN                : out   std_logic_vector(3 downto 0);                     -- arlen
			h2f_ARSIZE               : out   std_logic_vector(2 downto 0);                     -- arsize
			h2f_ARBURST              : out   std_logic_vector(1 downto 0);                     -- arburst
			h2f_ARLOCK               : out   std_logic_vector(1 downto 0);                     -- arlock
			h2f_ARCACHE              : out   std_logic_vector(3 downto 0);                     -- arcache
			h2f_ARPROT               : out   std_logic_vector(2 downto 0);                     -- arprot
			h2f_ARVALID              : out   std_logic;                                        -- arvalid
			h2f_ARREADY              : in    std_logic                     := 'X';             -- arready
			h2f_RID                  : in    std_logic_vector(11 downto 0) := (others => 'X'); -- rid
			h2f_RDATA                : in    std_logic_vector(63 downto 0) := (others => 'X'); -- rdata
			h2f_RRESP                : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			h2f_RLAST                : in    std_logic                     := 'X';             -- rlast
			h2f_RVALID               : in    std_logic                     := 'X';             -- rvalid
			h2f_RREADY               : out   std_logic;                                        -- rready
			h2f_lw_axi_clk           : in    std_logic                     := 'X';             -- clk
			h2f_lw_AWID              : out   std_logic_vector(11 downto 0);                    -- awid
			h2f_lw_AWADDR            : out   std_logic_vector(20 downto 0);                    -- awaddr
			h2f_lw_AWLEN             : out   std_logic_vector(3 downto 0);                     -- awlen
			h2f_lw_AWSIZE            : out   std_logic_vector(2 downto 0);                     -- awsize
			h2f_lw_AWBURST           : out   std_logic_vector(1 downto 0);                     -- awburst
			h2f_lw_AWLOCK            : out   std_logic_vector(1 downto 0);                     -- awlock
			h2f_lw_AWCACHE           : out   std_logic_vector(3 downto 0);                     -- awcache
			h2f_lw_AWPROT            : out   std_logic_vector(2 downto 0);                     -- awprot
			h2f_lw_AWVALID           : out   std_logic;                                        -- awvalid
			h2f_lw_AWREADY           : in    std_logic                     := 'X';             -- awready
			h2f_lw_WID               : out   std_logic_vector(11 downto 0);                    -- wid
			h2f_lw_WDATA             : out   std_logic_vector(31 downto 0);                    -- wdata
			h2f_lw_WSTRB             : out   std_logic_vector(3 downto 0);                     -- wstrb
			h2f_lw_WLAST             : out   std_logic;                                        -- wlast
			h2f_lw_WVALID            : out   std_logic;                                        -- wvalid
			h2f_lw_WREADY            : in    std_logic                     := 'X';             -- wready
			h2f_lw_BID               : in    std_logic_vector(11 downto 0) := (others => 'X'); -- bid
			h2f_lw_BRESP             : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			h2f_lw_BVALID            : in    std_logic                     := 'X';             -- bvalid
			h2f_lw_BREADY            : out   std_logic;                                        -- bready
			h2f_lw_ARID              : out   std_logic_vector(11 downto 0);                    -- arid
			h2f_lw_ARADDR            : out   std_logic_vector(20 downto 0);                    -- araddr
			h2f_lw_ARLEN             : out   std_logic_vector(3 downto 0);                     -- arlen
			h2f_lw_ARSIZE            : out   std_logic_vector(2 downto 0);                     -- arsize
			h2f_lw_ARBURST           : out   std_logic_vector(1 downto 0);                     -- arburst
			h2f_lw_ARLOCK            : out   std_logic_vector(1 downto 0);                     -- arlock
			h2f_lw_ARCACHE           : out   std_logic_vector(3 downto 0);                     -- arcache
			h2f_lw_ARPROT            : out   std_logic_vector(2 downto 0);                     -- arprot
			h2f_lw_ARVALID           : out   std_logic;                                        -- arvalid
			h2f_lw_ARREADY           : in    std_logic                     := 'X';             -- arready
			h2f_lw_RID               : in    std_logic_vector(11 downto 0) := (others => 'X'); -- rid
			h2f_lw_RDATA             : in    std_logic_vector(31 downto 0) := (others => 'X'); -- rdata
			h2f_lw_RRESP             : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			h2f_lw_RLAST             : in    std_logic                     := 'X';             -- rlast
			h2f_lw_RVALID            : in    std_logic                     := 'X';             -- rvalid
			h2f_lw_RREADY            : out   std_logic;                                        -- rready
			f2h_irq_p0               : in    std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			f2h_irq_p1               : in    std_logic_vector(31 downto 0) := (others => 'X')  -- irq
		);
	end component fluid_board_soc_hps_0;

	component fluid_board_soc_sysid is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component fluid_board_soc_sysid;

	component fluid_board_soc_pll_0 is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component fluid_board_soc_pll_0;

	component fluid_board_soc_sld_hub_controller_system_0 is
		generic (
			ENABLE_JTAG_IO_SELECTION : integer := 0
		);
		port (
			clk_clk          : in  std_logic                     := 'X';             -- clk
			reset_reset      : in  std_logic                     := 'X';             -- reset
			s0_waitrequest   : out std_logic;                                        -- waitrequest
			s0_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			s0_readdatavalid : out std_logic;                                        -- readdatavalid
			s0_burstcount    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			s0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			s0_address       : in  std_logic_vector(6 downto 0)  := (others => 'X'); -- address
			s0_write         : in  std_logic                     := 'X';             -- write
			s0_read          : in  std_logic                     := 'X';             -- read
			s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			s0_debugaccess   : in  std_logic                     := 'X'              -- debugaccess
		);
	end component fluid_board_soc_sld_hub_controller_system_0;

	component fluid_board_soc_nios2_qsys_0 is
		port (
			clk                                   : in  std_logic                     := 'X';             -- clk
			reset_n                               : in  std_logic                     := 'X';             -- reset_n
			reset_req                             : in  std_logic                     := 'X';             -- reset_req
			d_address                             : out std_logic_vector(18 downto 0);                    -- address
			d_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                                : out std_logic;                                        -- read
			d_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_write                               : out std_logic;                                        -- write
			d_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_debug_module_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                             : out std_logic_vector(16 downto 0);                    -- address
			i_read                                : out std_logic;                                        -- read
			i_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                       : in  std_logic                     := 'X';             -- readdatavalid
			d_irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			jtag_debug_module_resetrequest        : out std_logic;                                        -- reset
			jtag_debug_module_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			jtag_debug_module_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_debug_module_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			jtag_debug_module_read                : in  std_logic                     := 'X';             -- read
			jtag_debug_module_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_debug_module_waitrequest         : out std_logic;                                        -- waitrequest
			jtag_debug_module_write               : in  std_logic                     := 'X';             -- write
			jtag_debug_module_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			no_ci_readra                          : out std_logic;                                        -- readra
			cpu_resetrequest                      : in  std_logic                     := 'X';             -- export
			cpu_resettaken                        : out std_logic                                         -- export
		);
	end component fluid_board_soc_nios2_qsys_0;

	component fluid_board_soc_timer_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component fluid_board_soc_timer_0;

	component avalon_spi_AMC7891 is
		port (
			csi_clock_clk      : in  std_logic                     := 'X';             -- clk
			csi_clock_reset_n  : in  std_logic                     := 'X';             -- reset_n
			avs_s1_writedata   : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			avs_s1_read        : in  std_logic                     := 'X';             -- read
			avs_s1_write       : in  std_logic                     := 'X';             -- write
			avs_s1_address     : in  std_logic_vector(6 downto 0)  := (others => 'X'); -- address
			avs_s1_waitrequest : out std_logic;                                        -- waitrequest
			avs_s1_readdata    : out std_logic_vector(15 downto 0);                    -- readdata
			coe_s1_sclk        : out std_logic;                                        -- sclk
			coe_s1_cs_n        : out std_logic;                                        -- cs_n
			coe_s1_sdio        : out std_logic;                                        -- sdio
			coe_s1_sdo         : in  std_logic                     := 'X'              -- sdo
		);
	end component avalon_spi_AMC7891;

	component i2c_opencores is
		port (
			wb_adr_i   : in    std_logic_vector(2 downto 0) := (others => 'X'); -- address
			wb_dat_i   : in    std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			wb_dat_o   : out   std_logic_vector(7 downto 0);                    -- readdata
			wb_we_i    : in    std_logic                    := 'X';             -- write
			wb_stb_i   : in    std_logic                    := 'X';             -- chipselect
			wb_ack_o   : out   std_logic;                                       -- waitrequest_n
			scl_pad_io : inout std_logic                    := 'X';             -- scl
			sda_pad_io : inout std_logic                    := 'X';             -- sda
			wb_clk_i   : in    std_logic                    := 'X';             -- clk
			wb_rst_i   : in    std_logic                    := 'X';             -- reset
			wb_inta_o  : out   std_logic                                        -- irq
		);
	end component i2c_opencores;

	component fluid_board_soc_onchip_memory_nios_cpu is
		port (
			address     : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			clken       : in  std_logic                     := 'X';             -- clken
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			address2    : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			chipselect2 : in  std_logic                     := 'X';             -- chipselect
			clken2      : in  std_logic                     := 'X';             -- clken
			write2      : in  std_logic                     := 'X';             -- write
			readdata2   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata2  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable2 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			clk         : in  std_logic                     := 'X';             -- clk
			reset       : in  std_logic                     := 'X';             -- reset
			reset_req   : in  std_logic                     := 'X'              -- reset_req
		);
	end component fluid_board_soc_onchip_memory_nios_cpu;

	component fluid_board_soc_pio_input is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component fluid_board_soc_pio_input;

	component fluid_board_soc_pio_output is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component fluid_board_soc_pio_output;

	component fluid_board_soc_onchip_memory_nios_arm is
		port (
			address     : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			clken       : in  std_logic                     := 'X';             -- clken
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(15 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			byteenable  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			address2    : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			chipselect2 : in  std_logic                     := 'X';             -- chipselect
			clken2      : in  std_logic                     := 'X';             -- clken
			write2      : in  std_logic                     := 'X';             -- write
			readdata2   : out std_logic_vector(15 downto 0);                    -- readdata
			writedata2  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			byteenable2 : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			clk         : in  std_logic                     := 'X';             -- clk
			reset       : in  std_logic                     := 'X';             -- reset
			reset_req   : in  std_logic                     := 'X'              -- reset_req
		);
	end component fluid_board_soc_onchip_memory_nios_arm;

	component fluid_board_soc_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component fluid_board_soc_jtag_uart;

	component fluid_board_soc_fpga_only_master is
		port (
			clk_clk              : in  std_logic                     := 'X';             -- clk
			clk_reset_reset      : in  std_logic                     := 'X';             -- reset
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			master_read          : out std_logic;                                        -- read
			master_write         : out std_logic;                                        -- write
			master_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			master_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			master_reset_reset   : out std_logic                                         -- reset
		);
	end component fluid_board_soc_fpga_only_master;

	component fluid_board_soc_pio_reset_nios is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic                                         -- export
		);
	end component fluid_board_soc_pio_reset_nios;

	component fluid_board_soc_mm_interconnect_0 is
		port (
			hps_0_h2f_lw_axi_master_awid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- awid
			hps_0_h2f_lw_axi_master_awaddr                                      : in  std_logic_vector(20 downto 0) := (others => 'X'); -- awaddr
			hps_0_h2f_lw_axi_master_awlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awlen
			hps_0_h2f_lw_axi_master_awsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			hps_0_h2f_lw_axi_master_awburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awburst
			hps_0_h2f_lw_axi_master_awlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awlock
			hps_0_h2f_lw_axi_master_awcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awcache
			hps_0_h2f_lw_axi_master_awprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			hps_0_h2f_lw_axi_master_awvalid                                     : in  std_logic                     := 'X';             -- awvalid
			hps_0_h2f_lw_axi_master_awready                                     : out std_logic;                                        -- awready
			hps_0_h2f_lw_axi_master_wid                                         : in  std_logic_vector(11 downto 0) := (others => 'X'); -- wid
			hps_0_h2f_lw_axi_master_wdata                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wdata
			hps_0_h2f_lw_axi_master_wstrb                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- wstrb
			hps_0_h2f_lw_axi_master_wlast                                       : in  std_logic                     := 'X';             -- wlast
			hps_0_h2f_lw_axi_master_wvalid                                      : in  std_logic                     := 'X';             -- wvalid
			hps_0_h2f_lw_axi_master_wready                                      : out std_logic;                                        -- wready
			hps_0_h2f_lw_axi_master_bid                                         : out std_logic_vector(11 downto 0);                    -- bid
			hps_0_h2f_lw_axi_master_bresp                                       : out std_logic_vector(1 downto 0);                     -- bresp
			hps_0_h2f_lw_axi_master_bvalid                                      : out std_logic;                                        -- bvalid
			hps_0_h2f_lw_axi_master_bready                                      : in  std_logic                     := 'X';             -- bready
			hps_0_h2f_lw_axi_master_arid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- arid
			hps_0_h2f_lw_axi_master_araddr                                      : in  std_logic_vector(20 downto 0) := (others => 'X'); -- araddr
			hps_0_h2f_lw_axi_master_arlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arlen
			hps_0_h2f_lw_axi_master_arsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			hps_0_h2f_lw_axi_master_arburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arburst
			hps_0_h2f_lw_axi_master_arlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arlock
			hps_0_h2f_lw_axi_master_arcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arcache
			hps_0_h2f_lw_axi_master_arprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			hps_0_h2f_lw_axi_master_arvalid                                     : in  std_logic                     := 'X';             -- arvalid
			hps_0_h2f_lw_axi_master_arready                                     : out std_logic;                                        -- arready
			hps_0_h2f_lw_axi_master_rid                                         : out std_logic_vector(11 downto 0);                    -- rid
			hps_0_h2f_lw_axi_master_rdata                                       : out std_logic_vector(31 downto 0);                    -- rdata
			hps_0_h2f_lw_axi_master_rresp                                       : out std_logic_vector(1 downto 0);                     -- rresp
			hps_0_h2f_lw_axi_master_rlast                                       : out std_logic;                                        -- rlast
			hps_0_h2f_lw_axi_master_rvalid                                      : out std_logic;                                        -- rvalid
			hps_0_h2f_lw_axi_master_rready                                      : in  std_logic                     := 'X';             -- rready
			clk_i_clk_clk                                                       : in  std_logic                     := 'X';             -- clk
			fpga_only_master_clk_reset_reset_bridge_in_reset_reset              : in  std_logic                     := 'X';             -- reset
			hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			nios2_qsys_0_reset_n_reset_bridge_in_reset_reset                    : in  std_logic                     := 'X';             -- reset
			sysid_reset_reset_bridge_in_reset_reset                             : in  std_logic                     := 'X';             -- reset
			fpga_only_master_master_address                                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			fpga_only_master_master_waitrequest                                 : out std_logic;                                        -- waitrequest
			fpga_only_master_master_byteenable                                  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			fpga_only_master_master_read                                        : in  std_logic                     := 'X';             -- read
			fpga_only_master_master_readdata                                    : out std_logic_vector(31 downto 0);                    -- readdata
			fpga_only_master_master_readdatavalid                               : out std_logic;                                        -- readdatavalid
			fpga_only_master_master_write                                       : in  std_logic                     := 'X';             -- write
			fpga_only_master_master_writedata                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_qsys_0_data_master_address                                    : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address
			nios2_qsys_0_data_master_waitrequest                                : out std_logic;                                        -- waitrequest
			nios2_qsys_0_data_master_byteenable                                 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_qsys_0_data_master_read                                       : in  std_logic                     := 'X';             -- read
			nios2_qsys_0_data_master_readdata                                   : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_qsys_0_data_master_write                                      : in  std_logic                     := 'X';             -- write
			nios2_qsys_0_data_master_writedata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_qsys_0_data_master_debugaccess                                : in  std_logic                     := 'X';             -- debugaccess
			nios2_qsys_0_instruction_master_address                             : in  std_logic_vector(16 downto 0) := (others => 'X'); -- address
			nios2_qsys_0_instruction_master_waitrequest                         : out std_logic;                                        -- waitrequest
			nios2_qsys_0_instruction_master_read                                : in  std_logic                     := 'X';             -- read
			nios2_qsys_0_instruction_master_readdata                            : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_qsys_0_instruction_master_readdatavalid                       : out std_logic;                                        -- readdatavalid
			avalon_spi_AMC7891_0_s1_address                                     : out std_logic_vector(6 downto 0);                     -- address
			avalon_spi_AMC7891_0_s1_write                                       : out std_logic;                                        -- write
			avalon_spi_AMC7891_0_s1_read                                        : out std_logic;                                        -- read
			avalon_spi_AMC7891_0_s1_readdata                                    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			avalon_spi_AMC7891_0_s1_writedata                                   : out std_logic_vector(15 downto 0);                    -- writedata
			avalon_spi_AMC7891_0_s1_waitrequest                                 : in  std_logic                     := 'X';             -- waitrequest
			avalon_spi_AMC7891_1_s1_address                                     : out std_logic_vector(6 downto 0);                     -- address
			avalon_spi_AMC7891_1_s1_write                                       : out std_logic;                                        -- write
			avalon_spi_AMC7891_1_s1_read                                        : out std_logic;                                        -- read
			avalon_spi_AMC7891_1_s1_readdata                                    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			avalon_spi_AMC7891_1_s1_writedata                                   : out std_logic_vector(15 downto 0);                    -- writedata
			avalon_spi_AMC7891_1_s1_waitrequest                                 : in  std_logic                     := 'X';             -- waitrequest
			i2c_master_d_avalon_slave_0_address                                 : out std_logic_vector(2 downto 0);                     -- address
			i2c_master_d_avalon_slave_0_write                                   : out std_logic;                                        -- write
			i2c_master_d_avalon_slave_0_readdata                                : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			i2c_master_d_avalon_slave_0_writedata                               : out std_logic_vector(7 downto 0);                     -- writedata
			i2c_master_d_avalon_slave_0_waitrequest                             : in  std_logic                     := 'X';             -- waitrequest
			i2c_master_d_avalon_slave_0_chipselect                              : out std_logic;                                        -- chipselect
			i2c_master_f_avalon_slave_0_address                                 : out std_logic_vector(2 downto 0);                     -- address
			i2c_master_f_avalon_slave_0_write                                   : out std_logic;                                        -- write
			i2c_master_f_avalon_slave_0_readdata                                : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			i2c_master_f_avalon_slave_0_writedata                               : out std_logic_vector(7 downto 0);                     -- writedata
			i2c_master_f_avalon_slave_0_waitrequest                             : in  std_logic                     := 'X';             -- waitrequest
			i2c_master_f_avalon_slave_0_chipselect                              : out std_logic;                                        -- chipselect
			i2c_master_is1_avalon_slave_0_address                               : out std_logic_vector(2 downto 0);                     -- address
			i2c_master_is1_avalon_slave_0_write                                 : out std_logic;                                        -- write
			i2c_master_is1_avalon_slave_0_readdata                              : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			i2c_master_is1_avalon_slave_0_writedata                             : out std_logic_vector(7 downto 0);                     -- writedata
			i2c_master_is1_avalon_slave_0_waitrequest                           : in  std_logic                     := 'X';             -- waitrequest
			i2c_master_is1_avalon_slave_0_chipselect                            : out std_logic;                                        -- chipselect
			i2c_master_is2_avalon_slave_0_address                               : out std_logic_vector(2 downto 0);                     -- address
			i2c_master_is2_avalon_slave_0_write                                 : out std_logic;                                        -- write
			i2c_master_is2_avalon_slave_0_readdata                              : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			i2c_master_is2_avalon_slave_0_writedata                             : out std_logic_vector(7 downto 0);                     -- writedata
			i2c_master_is2_avalon_slave_0_waitrequest                           : in  std_logic                     := 'X';             -- waitrequest
			i2c_master_is2_avalon_slave_0_chipselect                            : out std_logic;                                        -- chipselect
			i2c_master_is3_avalon_slave_0_address                               : out std_logic_vector(2 downto 0);                     -- address
			i2c_master_is3_avalon_slave_0_write                                 : out std_logic;                                        -- write
			i2c_master_is3_avalon_slave_0_readdata                              : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			i2c_master_is3_avalon_slave_0_writedata                             : out std_logic_vector(7 downto 0);                     -- writedata
			i2c_master_is3_avalon_slave_0_waitrequest                           : in  std_logic                     := 'X';             -- waitrequest
			i2c_master_is3_avalon_slave_0_chipselect                            : out std_logic;                                        -- chipselect
			i2c_master_is4_avalon_slave_0_address                               : out std_logic_vector(2 downto 0);                     -- address
			i2c_master_is4_avalon_slave_0_write                                 : out std_logic;                                        -- write
			i2c_master_is4_avalon_slave_0_readdata                              : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			i2c_master_is4_avalon_slave_0_writedata                             : out std_logic_vector(7 downto 0);                     -- writedata
			i2c_master_is4_avalon_slave_0_waitrequest                           : in  std_logic                     := 'X';             -- waitrequest
			i2c_master_is4_avalon_slave_0_chipselect                            : out std_logic;                                        -- chipselect
			i2c_master_p_avalon_slave_0_address                                 : out std_logic_vector(2 downto 0);                     -- address
			i2c_master_p_avalon_slave_0_write                                   : out std_logic;                                        -- write
			i2c_master_p_avalon_slave_0_readdata                                : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			i2c_master_p_avalon_slave_0_writedata                               : out std_logic_vector(7 downto 0);                     -- writedata
			i2c_master_p_avalon_slave_0_waitrequest                             : in  std_logic                     := 'X';             -- waitrequest
			i2c_master_p_avalon_slave_0_chipselect                              : out std_logic;                                        -- chipselect
			jtag_uart_avalon_jtag_slave_address                                 : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write                                   : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read                                    : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest                             : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                              : out std_logic;                                        -- chipselect
			nios2_qsys_0_jtag_debug_module_address                              : out std_logic_vector(8 downto 0);                     -- address
			nios2_qsys_0_jtag_debug_module_write                                : out std_logic;                                        -- write
			nios2_qsys_0_jtag_debug_module_read                                 : out std_logic;                                        -- read
			nios2_qsys_0_jtag_debug_module_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_qsys_0_jtag_debug_module_writedata                            : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_qsys_0_jtag_debug_module_byteenable                           : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_qsys_0_jtag_debug_module_waitrequest                          : in  std_logic                     := 'X';             -- waitrequest
			nios2_qsys_0_jtag_debug_module_debugaccess                          : out std_logic;                                        -- debugaccess
			onchip_memory_nios_arm_s1_address                                   : out std_logic_vector(14 downto 0);                    -- address
			onchip_memory_nios_arm_s1_write                                     : out std_logic;                                        -- write
			onchip_memory_nios_arm_s1_readdata                                  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			onchip_memory_nios_arm_s1_writedata                                 : out std_logic_vector(15 downto 0);                    -- writedata
			onchip_memory_nios_arm_s1_byteenable                                : out std_logic_vector(1 downto 0);                     -- byteenable
			onchip_memory_nios_arm_s1_chipselect                                : out std_logic;                                        -- chipselect
			onchip_memory_nios_arm_s1_clken                                     : out std_logic;                                        -- clken
			onchip_memory_nios_cpu_s1_address                                   : out std_logic_vector(13 downto 0);                    -- address
			onchip_memory_nios_cpu_s1_write                                     : out std_logic;                                        -- write
			onchip_memory_nios_cpu_s1_readdata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory_nios_cpu_s1_writedata                                 : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory_nios_cpu_s1_byteenable                                : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory_nios_cpu_s1_chipselect                                : out std_logic;                                        -- chipselect
			onchip_memory_nios_cpu_s1_clken                                     : out std_logic;                                        -- clken
			pio_input_s1_address                                                : out std_logic_vector(1 downto 0);                     -- address
			pio_input_s1_write                                                  : out std_logic;                                        -- write
			pio_input_s1_readdata                                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_input_s1_writedata                                              : out std_logic_vector(31 downto 0);                    -- writedata
			pio_input_s1_chipselect                                             : out std_logic;                                        -- chipselect
			pio_output_s1_address                                               : out std_logic_vector(2 downto 0);                     -- address
			pio_output_s1_write                                                 : out std_logic;                                        -- write
			pio_output_s1_readdata                                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_output_s1_writedata                                             : out std_logic_vector(31 downto 0);                    -- writedata
			pio_output_s1_chipselect                                            : out std_logic;                                        -- chipselect
			pio_reset_nios_s1_address                                           : out std_logic_vector(1 downto 0);                     -- address
			pio_reset_nios_s1_write                                             : out std_logic;                                        -- write
			pio_reset_nios_s1_readdata                                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_reset_nios_s1_writedata                                         : out std_logic_vector(31 downto 0);                    -- writedata
			pio_reset_nios_s1_chipselect                                        : out std_logic;                                        -- chipselect
			sysid_control_slave_address                                         : out std_logic_vector(0 downto 0);                     -- address
			sysid_control_slave_readdata                                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			timer_0_s1_address                                                  : out std_logic_vector(2 downto 0);                     -- address
			timer_0_s1_write                                                    : out std_logic;                                        -- write
			timer_0_s1_readdata                                                 : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_0_s1_writedata                                                : out std_logic_vector(15 downto 0);                    -- writedata
			timer_0_s1_chipselect                                               : out std_logic;                                        -- chipselect
			timer_1_s1_address                                                  : out std_logic_vector(2 downto 0);                     -- address
			timer_1_s1_write                                                    : out std_logic;                                        -- write
			timer_1_s1_readdata                                                 : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_1_s1_writedata                                                : out std_logic_vector(15 downto 0);                    -- writedata
			timer_1_s1_chipselect                                               : out std_logic                                         -- chipselect
		);
	end component fluid_board_soc_mm_interconnect_0;

	component fluid_board_soc_mm_interconnect_1 is
		port (
			hps_0_h2f_axi_master_awid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- awid
			hps_0_h2f_axi_master_awaddr                                      : in  std_logic_vector(29 downto 0) := (others => 'X'); -- awaddr
			hps_0_h2f_axi_master_awlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awlen
			hps_0_h2f_axi_master_awsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			hps_0_h2f_axi_master_awburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awburst
			hps_0_h2f_axi_master_awlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awlock
			hps_0_h2f_axi_master_awcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awcache
			hps_0_h2f_axi_master_awprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			hps_0_h2f_axi_master_awvalid                                     : in  std_logic                     := 'X';             -- awvalid
			hps_0_h2f_axi_master_awready                                     : out std_logic;                                        -- awready
			hps_0_h2f_axi_master_wid                                         : in  std_logic_vector(11 downto 0) := (others => 'X'); -- wid
			hps_0_h2f_axi_master_wdata                                       : in  std_logic_vector(63 downto 0) := (others => 'X'); -- wdata
			hps_0_h2f_axi_master_wstrb                                       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wstrb
			hps_0_h2f_axi_master_wlast                                       : in  std_logic                     := 'X';             -- wlast
			hps_0_h2f_axi_master_wvalid                                      : in  std_logic                     := 'X';             -- wvalid
			hps_0_h2f_axi_master_wready                                      : out std_logic;                                        -- wready
			hps_0_h2f_axi_master_bid                                         : out std_logic_vector(11 downto 0);                    -- bid
			hps_0_h2f_axi_master_bresp                                       : out std_logic_vector(1 downto 0);                     -- bresp
			hps_0_h2f_axi_master_bvalid                                      : out std_logic;                                        -- bvalid
			hps_0_h2f_axi_master_bready                                      : in  std_logic                     := 'X';             -- bready
			hps_0_h2f_axi_master_arid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- arid
			hps_0_h2f_axi_master_araddr                                      : in  std_logic_vector(29 downto 0) := (others => 'X'); -- araddr
			hps_0_h2f_axi_master_arlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arlen
			hps_0_h2f_axi_master_arsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			hps_0_h2f_axi_master_arburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arburst
			hps_0_h2f_axi_master_arlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arlock
			hps_0_h2f_axi_master_arcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arcache
			hps_0_h2f_axi_master_arprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			hps_0_h2f_axi_master_arvalid                                     : in  std_logic                     := 'X';             -- arvalid
			hps_0_h2f_axi_master_arready                                     : out std_logic;                                        -- arready
			hps_0_h2f_axi_master_rid                                         : out std_logic_vector(11 downto 0);                    -- rid
			hps_0_h2f_axi_master_rdata                                       : out std_logic_vector(63 downto 0);                    -- rdata
			hps_0_h2f_axi_master_rresp                                       : out std_logic_vector(1 downto 0);                     -- rresp
			hps_0_h2f_axi_master_rlast                                       : out std_logic;                                        -- rlast
			hps_0_h2f_axi_master_rvalid                                      : out std_logic;                                        -- rvalid
			hps_0_h2f_axi_master_rready                                      : in  std_logic                     := 'X';             -- rready
			clk_i_clk_clk                                                    : in  std_logic                     := 'X';             -- clk
			hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			sld_hub_controller_system_0_reset_reset_bridge_in_reset_reset    : in  std_logic                     := 'X';             -- reset
			onchip_memory_nios_arm_s2_address                                : out std_logic_vector(14 downto 0);                    -- address
			onchip_memory_nios_arm_s2_write                                  : out std_logic;                                        -- write
			onchip_memory_nios_arm_s2_readdata                               : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			onchip_memory_nios_arm_s2_writedata                              : out std_logic_vector(15 downto 0);                    -- writedata
			onchip_memory_nios_arm_s2_byteenable                             : out std_logic_vector(1 downto 0);                     -- byteenable
			onchip_memory_nios_arm_s2_chipselect                             : out std_logic;                                        -- chipselect
			onchip_memory_nios_arm_s2_clken                                  : out std_logic;                                        -- clken
			onchip_memory_nios_cpu_s2_address                                : out std_logic_vector(13 downto 0);                    -- address
			onchip_memory_nios_cpu_s2_write                                  : out std_logic;                                        -- write
			onchip_memory_nios_cpu_s2_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory_nios_cpu_s2_writedata                              : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory_nios_cpu_s2_byteenable                             : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory_nios_cpu_s2_chipselect                             : out std_logic;                                        -- chipselect
			onchip_memory_nios_cpu_s2_clken                                  : out std_logic;                                        -- clken
			sld_hub_controller_system_0_s0_address                           : out std_logic_vector(6 downto 0);                     -- address
			sld_hub_controller_system_0_s0_write                             : out std_logic;                                        -- write
			sld_hub_controller_system_0_s0_read                              : out std_logic;                                        -- read
			sld_hub_controller_system_0_s0_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sld_hub_controller_system_0_s0_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			sld_hub_controller_system_0_s0_burstcount                        : out std_logic_vector(0 downto 0);                     -- burstcount
			sld_hub_controller_system_0_s0_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			sld_hub_controller_system_0_s0_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			sld_hub_controller_system_0_s0_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			sld_hub_controller_system_0_s0_debugaccess                       : out std_logic                                         -- debugaccess
		);
	end component fluid_board_soc_mm_interconnect_1;

	component fluid_board_soc_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component fluid_board_soc_irq_mapper;

	component fluid_board_soc_irq_mapper_001 is
		port (
			clk        : in  std_logic                     := 'X'; -- clk
			reset      : in  std_logic                     := 'X'; -- reset
			sender_irq : out std_logic_vector(31 downto 0)         -- irq
		);
	end component fluid_board_soc_irq_mapper_001;

	component fluid_board_soc_irq_mapper_002 is
		port (
			clk            : in  std_logic                     := 'X'; -- clk
			reset          : in  std_logic                     := 'X'; -- reset
			receiver0_irq  : in  std_logic                     := 'X'; -- irq
			receiver1_irq  : in  std_logic                     := 'X'; -- irq
			receiver2_irq  : in  std_logic                     := 'X'; -- irq
			receiver3_irq  : in  std_logic                     := 'X'; -- irq
			receiver4_irq  : in  std_logic                     := 'X'; -- irq
			receiver5_irq  : in  std_logic                     := 'X'; -- irq
			receiver6_irq  : in  std_logic                     := 'X'; -- irq
			receiver7_irq  : in  std_logic                     := 'X'; -- irq
			receiver8_irq  : in  std_logic                     := 'X'; -- irq
			receiver9_irq  : in  std_logic                     := 'X'; -- irq
			receiver10_irq : in  std_logic                     := 'X'; -- irq
			sender_irq     : out std_logic_vector(31 downto 0)         -- irq
		);
	end component fluid_board_soc_irq_mapper_002;

	component fluid_board_soc_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component fluid_board_soc_rst_controller;

	component fluid_board_soc_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component fluid_board_soc_rst_controller_001;

	component fluid_board_soc_rst_controller_002 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component fluid_board_soc_rst_controller_002;

	signal pll_0_outclk0_clk                                              : std_logic;                     -- pll_0:outclk_0 -> [pll_0_sys_clk_clk, avalon_spi_AMC7891_0:csi_clock_clk, avalon_spi_AMC7891_1:csi_clock_clk, fpga_only_master:clk_clk, hps_0:h2f_axi_clk, hps_0:h2f_lw_axi_clk, i2c_master_d:wb_clk_i, i2c_master_f:wb_clk_i, i2c_master_is1:wb_clk_i, i2c_master_is2:wb_clk_i, i2c_master_is3:wb_clk_i, i2c_master_is4:wb_clk_i, i2c_master_p:wb_clk_i, irq_mapper_002:clk, jtag_uart:clk, mm_interconnect_0:clk_i_clk_clk, mm_interconnect_1:clk_i_clk_clk, nios2_qsys_0:clk, onchip_memory_nios_arm:clk, onchip_memory_nios_cpu:clk, pio_input:clk, pio_output:clk, pio_reset_nios:clk, rst_controller:clk, rst_controller_001:clk, rst_controller_002:clk, sld_hub_controller_system_0:clk_clk, sysid:clock, timer_0:clk, timer_1:clk]
	signal hps_0_h2f_lw_axi_master_awvalid                                : std_logic;                     -- hps_0:h2f_lw_AWVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awvalid
	signal hps_0_h2f_lw_axi_master_arsize                                 : std_logic_vector(2 downto 0);  -- hps_0:h2f_lw_ARSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arsize
	signal hps_0_h2f_lw_axi_master_arlock                                 : std_logic_vector(1 downto 0);  -- hps_0:h2f_lw_ARLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlock
	signal hps_0_h2f_lw_axi_master_awcache                                : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_AWCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awcache
	signal hps_0_h2f_lw_axi_master_arready                                : std_logic;                     -- mm_interconnect_0:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	signal hps_0_h2f_lw_axi_master_arid                                   : std_logic_vector(11 downto 0); -- hps_0:h2f_lw_ARID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arid
	signal hps_0_h2f_lw_axi_master_rready                                 : std_logic;                     -- hps_0:h2f_lw_RREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_rready
	signal hps_0_h2f_lw_axi_master_bready                                 : std_logic;                     -- hps_0:h2f_lw_BREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_bready
	signal hps_0_h2f_lw_axi_master_awsize                                 : std_logic_vector(2 downto 0);  -- hps_0:h2f_lw_AWSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awsize
	signal hps_0_h2f_lw_axi_master_awprot                                 : std_logic_vector(2 downto 0);  -- hps_0:h2f_lw_AWPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awprot
	signal hps_0_h2f_lw_axi_master_arvalid                                : std_logic;                     -- hps_0:h2f_lw_ARVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arvalid
	signal hps_0_h2f_lw_axi_master_arprot                                 : std_logic_vector(2 downto 0);  -- hps_0:h2f_lw_ARPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arprot
	signal hps_0_h2f_lw_axi_master_bid                                    : std_logic_vector(11 downto 0); -- mm_interconnect_0:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	signal hps_0_h2f_lw_axi_master_arlen                                  : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_ARLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlen
	signal hps_0_h2f_lw_axi_master_awready                                : std_logic;                     -- mm_interconnect_0:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	signal hps_0_h2f_lw_axi_master_awid                                   : std_logic_vector(11 downto 0); -- hps_0:h2f_lw_AWID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awid
	signal hps_0_h2f_lw_axi_master_bvalid                                 : std_logic;                     -- mm_interconnect_0:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	signal hps_0_h2f_lw_axi_master_wid                                    : std_logic_vector(11 downto 0); -- hps_0:h2f_lw_WID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wid
	signal hps_0_h2f_lw_axi_master_awlock                                 : std_logic_vector(1 downto 0);  -- hps_0:h2f_lw_AWLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlock
	signal hps_0_h2f_lw_axi_master_awburst                                : std_logic_vector(1 downto 0);  -- hps_0:h2f_lw_AWBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awburst
	signal hps_0_h2f_lw_axi_master_bresp                                  : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	signal hps_0_h2f_lw_axi_master_wstrb                                  : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_WSTRB -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wstrb
	signal hps_0_h2f_lw_axi_master_rvalid                                 : std_logic;                     -- mm_interconnect_0:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	signal hps_0_h2f_lw_axi_master_wdata                                  : std_logic_vector(31 downto 0); -- hps_0:h2f_lw_WDATA -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wdata
	signal hps_0_h2f_lw_axi_master_wready                                 : std_logic;                     -- mm_interconnect_0:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	signal hps_0_h2f_lw_axi_master_arburst                                : std_logic_vector(1 downto 0);  -- hps_0:h2f_lw_ARBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arburst
	signal hps_0_h2f_lw_axi_master_rdata                                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	signal hps_0_h2f_lw_axi_master_araddr                                 : std_logic_vector(20 downto 0); -- hps_0:h2f_lw_ARADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_araddr
	signal hps_0_h2f_lw_axi_master_arcache                                : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_ARCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arcache
	signal hps_0_h2f_lw_axi_master_awlen                                  : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_AWLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlen
	signal hps_0_h2f_lw_axi_master_awaddr                                 : std_logic_vector(20 downto 0); -- hps_0:h2f_lw_AWADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awaddr
	signal hps_0_h2f_lw_axi_master_rid                                    : std_logic_vector(11 downto 0); -- mm_interconnect_0:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	signal hps_0_h2f_lw_axi_master_wvalid                                 : std_logic;                     -- hps_0:h2f_lw_WVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wvalid
	signal hps_0_h2f_lw_axi_master_rresp                                  : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	signal hps_0_h2f_lw_axi_master_wlast                                  : std_logic;                     -- hps_0:h2f_lw_WLAST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wlast
	signal hps_0_h2f_lw_axi_master_rlast                                  : std_logic;                     -- mm_interconnect_0:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	signal fpga_only_master_master_waitrequest                            : std_logic;                     -- mm_interconnect_0:fpga_only_master_master_waitrequest -> fpga_only_master:master_waitrequest
	signal fpga_only_master_master_writedata                              : std_logic_vector(31 downto 0); -- fpga_only_master:master_writedata -> mm_interconnect_0:fpga_only_master_master_writedata
	signal fpga_only_master_master_address                                : std_logic_vector(31 downto 0); -- fpga_only_master:master_address -> mm_interconnect_0:fpga_only_master_master_address
	signal fpga_only_master_master_write                                  : std_logic;                     -- fpga_only_master:master_write -> mm_interconnect_0:fpga_only_master_master_write
	signal fpga_only_master_master_read                                   : std_logic;                     -- fpga_only_master:master_read -> mm_interconnect_0:fpga_only_master_master_read
	signal fpga_only_master_master_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:fpga_only_master_master_readdata -> fpga_only_master:master_readdata
	signal fpga_only_master_master_byteenable                             : std_logic_vector(3 downto 0);  -- fpga_only_master:master_byteenable -> mm_interconnect_0:fpga_only_master_master_byteenable
	signal fpga_only_master_master_readdatavalid                          : std_logic;                     -- mm_interconnect_0:fpga_only_master_master_readdatavalid -> fpga_only_master:master_readdatavalid
	signal nios2_qsys_0_data_master_waitrequest                           : std_logic;                     -- mm_interconnect_0:nios2_qsys_0_data_master_waitrequest -> nios2_qsys_0:d_waitrequest
	signal nios2_qsys_0_data_master_writedata                             : std_logic_vector(31 downto 0); -- nios2_qsys_0:d_writedata -> mm_interconnect_0:nios2_qsys_0_data_master_writedata
	signal nios2_qsys_0_data_master_address                               : std_logic_vector(18 downto 0); -- nios2_qsys_0:d_address -> mm_interconnect_0:nios2_qsys_0_data_master_address
	signal nios2_qsys_0_data_master_write                                 : std_logic;                     -- nios2_qsys_0:d_write -> mm_interconnect_0:nios2_qsys_0_data_master_write
	signal nios2_qsys_0_data_master_read                                  : std_logic;                     -- nios2_qsys_0:d_read -> mm_interconnect_0:nios2_qsys_0_data_master_read
	signal nios2_qsys_0_data_master_readdata                              : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_qsys_0_data_master_readdata -> nios2_qsys_0:d_readdata
	signal nios2_qsys_0_data_master_debugaccess                           : std_logic;                     -- nios2_qsys_0:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_0_data_master_debugaccess
	signal nios2_qsys_0_data_master_byteenable                            : std_logic_vector(3 downto 0);  -- nios2_qsys_0:d_byteenable -> mm_interconnect_0:nios2_qsys_0_data_master_byteenable
	signal nios2_qsys_0_instruction_master_waitrequest                    : std_logic;                     -- mm_interconnect_0:nios2_qsys_0_instruction_master_waitrequest -> nios2_qsys_0:i_waitrequest
	signal nios2_qsys_0_instruction_master_address                        : std_logic_vector(16 downto 0); -- nios2_qsys_0:i_address -> mm_interconnect_0:nios2_qsys_0_instruction_master_address
	signal nios2_qsys_0_instruction_master_read                           : std_logic;                     -- nios2_qsys_0:i_read -> mm_interconnect_0:nios2_qsys_0_instruction_master_read
	signal nios2_qsys_0_instruction_master_readdata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_qsys_0_instruction_master_readdata -> nios2_qsys_0:i_readdata
	signal nios2_qsys_0_instruction_master_readdatavalid                  : std_logic;                     -- mm_interconnect_0:nios2_qsys_0_instruction_master_readdatavalid -> nios2_qsys_0:i_readdatavalid
	signal mm_interconnect_0_sysid_control_slave_address                  : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_control_slave_address -> sysid:address
	signal mm_interconnect_0_sysid_control_slave_readdata                 : std_logic_vector(31 downto 0); -- sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest      : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata        : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address          : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect       : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write            : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read             : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata         : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_0_pio_reset_nios_s1_writedata                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_reset_nios_s1_writedata -> pio_reset_nios:writedata
	signal mm_interconnect_0_pio_reset_nios_s1_address                    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_reset_nios_s1_address -> pio_reset_nios:address
	signal mm_interconnect_0_pio_reset_nios_s1_chipselect                 : std_logic;                     -- mm_interconnect_0:pio_reset_nios_s1_chipselect -> pio_reset_nios:chipselect
	signal mm_interconnect_0_pio_reset_nios_s1_write                      : std_logic;                     -- mm_interconnect_0:pio_reset_nios_s1_write -> mm_interconnect_0_pio_reset_nios_s1_write:in
	signal mm_interconnect_0_pio_reset_nios_s1_readdata                   : std_logic_vector(31 downto 0); -- pio_reset_nios:readdata -> mm_interconnect_0:pio_reset_nios_s1_readdata
	signal mm_interconnect_0_onchip_memory_nios_cpu_s1_writedata          : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory_nios_cpu_s1_writedata -> onchip_memory_nios_cpu:writedata
	signal mm_interconnect_0_onchip_memory_nios_cpu_s1_address            : std_logic_vector(13 downto 0); -- mm_interconnect_0:onchip_memory_nios_cpu_s1_address -> onchip_memory_nios_cpu:address
	signal mm_interconnect_0_onchip_memory_nios_cpu_s1_chipselect         : std_logic;                     -- mm_interconnect_0:onchip_memory_nios_cpu_s1_chipselect -> onchip_memory_nios_cpu:chipselect
	signal mm_interconnect_0_onchip_memory_nios_cpu_s1_clken              : std_logic;                     -- mm_interconnect_0:onchip_memory_nios_cpu_s1_clken -> onchip_memory_nios_cpu:clken
	signal mm_interconnect_0_onchip_memory_nios_cpu_s1_write              : std_logic;                     -- mm_interconnect_0:onchip_memory_nios_cpu_s1_write -> onchip_memory_nios_cpu:write
	signal mm_interconnect_0_onchip_memory_nios_cpu_s1_readdata           : std_logic_vector(31 downto 0); -- onchip_memory_nios_cpu:readdata -> mm_interconnect_0:onchip_memory_nios_cpu_s1_readdata
	signal mm_interconnect_0_onchip_memory_nios_cpu_s1_byteenable         : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory_nios_cpu_s1_byteenable -> onchip_memory_nios_cpu:byteenable
	signal mm_interconnect_0_onchip_memory_nios_arm_s1_writedata          : std_logic_vector(15 downto 0); -- mm_interconnect_0:onchip_memory_nios_arm_s1_writedata -> onchip_memory_nios_arm:writedata
	signal mm_interconnect_0_onchip_memory_nios_arm_s1_address            : std_logic_vector(14 downto 0); -- mm_interconnect_0:onchip_memory_nios_arm_s1_address -> onchip_memory_nios_arm:address
	signal mm_interconnect_0_onchip_memory_nios_arm_s1_chipselect         : std_logic;                     -- mm_interconnect_0:onchip_memory_nios_arm_s1_chipselect -> onchip_memory_nios_arm:chipselect
	signal mm_interconnect_0_onchip_memory_nios_arm_s1_clken              : std_logic;                     -- mm_interconnect_0:onchip_memory_nios_arm_s1_clken -> onchip_memory_nios_arm:clken
	signal mm_interconnect_0_onchip_memory_nios_arm_s1_write              : std_logic;                     -- mm_interconnect_0:onchip_memory_nios_arm_s1_write -> onchip_memory_nios_arm:write
	signal mm_interconnect_0_onchip_memory_nios_arm_s1_readdata           : std_logic_vector(15 downto 0); -- onchip_memory_nios_arm:readdata -> mm_interconnect_0:onchip_memory_nios_arm_s1_readdata
	signal mm_interconnect_0_onchip_memory_nios_arm_s1_byteenable         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:onchip_memory_nios_arm_s1_byteenable -> onchip_memory_nios_arm:byteenable
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest   : std_logic;                     -- nios2_qsys_0:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_waitrequest
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata     : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_qsys_0_jtag_debug_module_writedata -> nios2_qsys_0:jtag_debug_module_writedata
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address       : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_qsys_0_jtag_debug_module_address -> nios2_qsys_0:jtag_debug_module_address
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write         : std_logic;                     -- mm_interconnect_0:nios2_qsys_0_jtag_debug_module_write -> nios2_qsys_0:jtag_debug_module_write
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read          : std_logic;                     -- mm_interconnect_0:nios2_qsys_0_jtag_debug_module_read -> nios2_qsys_0:jtag_debug_module_read
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata      : std_logic_vector(31 downto 0); -- nios2_qsys_0:jtag_debug_module_readdata -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_readdata
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess   : std_logic;                     -- mm_interconnect_0:nios2_qsys_0_jtag_debug_module_debugaccess -> nios2_qsys_0:jtag_debug_module_debugaccess
	signal mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable    : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_qsys_0_jtag_debug_module_byteenable -> nios2_qsys_0:jtag_debug_module_byteenable
	signal mm_interconnect_0_timer_0_s1_writedata                         : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	signal mm_interconnect_0_timer_0_s1_address                           : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer_0_s1_address -> timer_0:address
	signal mm_interconnect_0_timer_0_s1_chipselect                        : std_logic;                     -- mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	signal mm_interconnect_0_timer_0_s1_write                             : std_logic;                     -- mm_interconnect_0:timer_0_s1_write -> mm_interconnect_0_timer_0_s1_write:in
	signal mm_interconnect_0_timer_0_s1_readdata                          : std_logic_vector(15 downto 0); -- timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	signal mm_interconnect_0_timer_1_s1_writedata                         : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_1_s1_writedata -> timer_1:writedata
	signal mm_interconnect_0_timer_1_s1_address                           : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer_1_s1_address -> timer_1:address
	signal mm_interconnect_0_timer_1_s1_chipselect                        : std_logic;                     -- mm_interconnect_0:timer_1_s1_chipselect -> timer_1:chipselect
	signal mm_interconnect_0_timer_1_s1_write                             : std_logic;                     -- mm_interconnect_0:timer_1_s1_write -> mm_interconnect_0_timer_1_s1_write:in
	signal mm_interconnect_0_timer_1_s1_readdata                          : std_logic_vector(15 downto 0); -- timer_1:readdata -> mm_interconnect_0:timer_1_s1_readdata
	signal mm_interconnect_0_avalon_spi_amc7891_0_s1_waitrequest          : std_logic;                     -- avalon_spi_AMC7891_0:avs_s1_waitrequest -> mm_interconnect_0:avalon_spi_AMC7891_0_s1_waitrequest
	signal mm_interconnect_0_avalon_spi_amc7891_0_s1_writedata            : std_logic_vector(15 downto 0); -- mm_interconnect_0:avalon_spi_AMC7891_0_s1_writedata -> avalon_spi_AMC7891_0:avs_s1_writedata
	signal mm_interconnect_0_avalon_spi_amc7891_0_s1_address              : std_logic_vector(6 downto 0);  -- mm_interconnect_0:avalon_spi_AMC7891_0_s1_address -> avalon_spi_AMC7891_0:avs_s1_address
	signal mm_interconnect_0_avalon_spi_amc7891_0_s1_write                : std_logic;                     -- mm_interconnect_0:avalon_spi_AMC7891_0_s1_write -> avalon_spi_AMC7891_0:avs_s1_write
	signal mm_interconnect_0_avalon_spi_amc7891_0_s1_read                 : std_logic;                     -- mm_interconnect_0:avalon_spi_AMC7891_0_s1_read -> avalon_spi_AMC7891_0:avs_s1_read
	signal mm_interconnect_0_avalon_spi_amc7891_0_s1_readdata             : std_logic_vector(15 downto 0); -- avalon_spi_AMC7891_0:avs_s1_readdata -> mm_interconnect_0:avalon_spi_AMC7891_0_s1_readdata
	signal mm_interconnect_0_avalon_spi_amc7891_1_s1_waitrequest          : std_logic;                     -- avalon_spi_AMC7891_1:avs_s1_waitrequest -> mm_interconnect_0:avalon_spi_AMC7891_1_s1_waitrequest
	signal mm_interconnect_0_avalon_spi_amc7891_1_s1_writedata            : std_logic_vector(15 downto 0); -- mm_interconnect_0:avalon_spi_AMC7891_1_s1_writedata -> avalon_spi_AMC7891_1:avs_s1_writedata
	signal mm_interconnect_0_avalon_spi_amc7891_1_s1_address              : std_logic_vector(6 downto 0);  -- mm_interconnect_0:avalon_spi_AMC7891_1_s1_address -> avalon_spi_AMC7891_1:avs_s1_address
	signal mm_interconnect_0_avalon_spi_amc7891_1_s1_write                : std_logic;                     -- mm_interconnect_0:avalon_spi_AMC7891_1_s1_write -> avalon_spi_AMC7891_1:avs_s1_write
	signal mm_interconnect_0_avalon_spi_amc7891_1_s1_read                 : std_logic;                     -- mm_interconnect_0:avalon_spi_AMC7891_1_s1_read -> avalon_spi_AMC7891_1:avs_s1_read
	signal mm_interconnect_0_avalon_spi_amc7891_1_s1_readdata             : std_logic_vector(15 downto 0); -- avalon_spi_AMC7891_1:avs_s1_readdata -> mm_interconnect_0:avalon_spi_AMC7891_1_s1_readdata
	signal i2c_master_is1_avalon_slave_0_waitrequest                      : std_logic;                     -- i2c_master_is1:wb_ack_o -> i2c_master_is1_avalon_slave_0_waitrequest:in
	signal mm_interconnect_0_i2c_master_is1_avalon_slave_0_writedata      : std_logic_vector(7 downto 0);  -- mm_interconnect_0:i2c_master_is1_avalon_slave_0_writedata -> i2c_master_is1:wb_dat_i
	signal mm_interconnect_0_i2c_master_is1_avalon_slave_0_address        : std_logic_vector(2 downto 0);  -- mm_interconnect_0:i2c_master_is1_avalon_slave_0_address -> i2c_master_is1:wb_adr_i
	signal mm_interconnect_0_i2c_master_is1_avalon_slave_0_chipselect     : std_logic;                     -- mm_interconnect_0:i2c_master_is1_avalon_slave_0_chipselect -> i2c_master_is1:wb_stb_i
	signal mm_interconnect_0_i2c_master_is1_avalon_slave_0_write          : std_logic;                     -- mm_interconnect_0:i2c_master_is1_avalon_slave_0_write -> i2c_master_is1:wb_we_i
	signal mm_interconnect_0_i2c_master_is1_avalon_slave_0_readdata       : std_logic_vector(7 downto 0);  -- i2c_master_is1:wb_dat_o -> mm_interconnect_0:i2c_master_is1_avalon_slave_0_readdata
	signal i2c_master_is2_avalon_slave_0_waitrequest                      : std_logic;                     -- i2c_master_is2:wb_ack_o -> i2c_master_is2_avalon_slave_0_waitrequest:in
	signal mm_interconnect_0_i2c_master_is2_avalon_slave_0_writedata      : std_logic_vector(7 downto 0);  -- mm_interconnect_0:i2c_master_is2_avalon_slave_0_writedata -> i2c_master_is2:wb_dat_i
	signal mm_interconnect_0_i2c_master_is2_avalon_slave_0_address        : std_logic_vector(2 downto 0);  -- mm_interconnect_0:i2c_master_is2_avalon_slave_0_address -> i2c_master_is2:wb_adr_i
	signal mm_interconnect_0_i2c_master_is2_avalon_slave_0_chipselect     : std_logic;                     -- mm_interconnect_0:i2c_master_is2_avalon_slave_0_chipselect -> i2c_master_is2:wb_stb_i
	signal mm_interconnect_0_i2c_master_is2_avalon_slave_0_write          : std_logic;                     -- mm_interconnect_0:i2c_master_is2_avalon_slave_0_write -> i2c_master_is2:wb_we_i
	signal mm_interconnect_0_i2c_master_is2_avalon_slave_0_readdata       : std_logic_vector(7 downto 0);  -- i2c_master_is2:wb_dat_o -> mm_interconnect_0:i2c_master_is2_avalon_slave_0_readdata
	signal i2c_master_is3_avalon_slave_0_waitrequest                      : std_logic;                     -- i2c_master_is3:wb_ack_o -> i2c_master_is3_avalon_slave_0_waitrequest:in
	signal mm_interconnect_0_i2c_master_is3_avalon_slave_0_writedata      : std_logic_vector(7 downto 0);  -- mm_interconnect_0:i2c_master_is3_avalon_slave_0_writedata -> i2c_master_is3:wb_dat_i
	signal mm_interconnect_0_i2c_master_is3_avalon_slave_0_address        : std_logic_vector(2 downto 0);  -- mm_interconnect_0:i2c_master_is3_avalon_slave_0_address -> i2c_master_is3:wb_adr_i
	signal mm_interconnect_0_i2c_master_is3_avalon_slave_0_chipselect     : std_logic;                     -- mm_interconnect_0:i2c_master_is3_avalon_slave_0_chipselect -> i2c_master_is3:wb_stb_i
	signal mm_interconnect_0_i2c_master_is3_avalon_slave_0_write          : std_logic;                     -- mm_interconnect_0:i2c_master_is3_avalon_slave_0_write -> i2c_master_is3:wb_we_i
	signal mm_interconnect_0_i2c_master_is3_avalon_slave_0_readdata       : std_logic_vector(7 downto 0);  -- i2c_master_is3:wb_dat_o -> mm_interconnect_0:i2c_master_is3_avalon_slave_0_readdata
	signal i2c_master_is4_avalon_slave_0_waitrequest                      : std_logic;                     -- i2c_master_is4:wb_ack_o -> i2c_master_is4_avalon_slave_0_waitrequest:in
	signal mm_interconnect_0_i2c_master_is4_avalon_slave_0_writedata      : std_logic_vector(7 downto 0);  -- mm_interconnect_0:i2c_master_is4_avalon_slave_0_writedata -> i2c_master_is4:wb_dat_i
	signal mm_interconnect_0_i2c_master_is4_avalon_slave_0_address        : std_logic_vector(2 downto 0);  -- mm_interconnect_0:i2c_master_is4_avalon_slave_0_address -> i2c_master_is4:wb_adr_i
	signal mm_interconnect_0_i2c_master_is4_avalon_slave_0_chipselect     : std_logic;                     -- mm_interconnect_0:i2c_master_is4_avalon_slave_0_chipselect -> i2c_master_is4:wb_stb_i
	signal mm_interconnect_0_i2c_master_is4_avalon_slave_0_write          : std_logic;                     -- mm_interconnect_0:i2c_master_is4_avalon_slave_0_write -> i2c_master_is4:wb_we_i
	signal mm_interconnect_0_i2c_master_is4_avalon_slave_0_readdata       : std_logic_vector(7 downto 0);  -- i2c_master_is4:wb_dat_o -> mm_interconnect_0:i2c_master_is4_avalon_slave_0_readdata
	signal mm_interconnect_0_pio_input_s1_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_input_s1_writedata -> pio_input:writedata
	signal mm_interconnect_0_pio_input_s1_address                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_input_s1_address -> pio_input:address
	signal mm_interconnect_0_pio_input_s1_chipselect                      : std_logic;                     -- mm_interconnect_0:pio_input_s1_chipselect -> pio_input:chipselect
	signal mm_interconnect_0_pio_input_s1_write                           : std_logic;                     -- mm_interconnect_0:pio_input_s1_write -> mm_interconnect_0_pio_input_s1_write:in
	signal mm_interconnect_0_pio_input_s1_readdata                        : std_logic_vector(31 downto 0); -- pio_input:readdata -> mm_interconnect_0:pio_input_s1_readdata
	signal mm_interconnect_0_pio_output_s1_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_output_s1_writedata -> pio_output:writedata
	signal mm_interconnect_0_pio_output_s1_address                        : std_logic_vector(2 downto 0);  -- mm_interconnect_0:pio_output_s1_address -> pio_output:address
	signal mm_interconnect_0_pio_output_s1_chipselect                     : std_logic;                     -- mm_interconnect_0:pio_output_s1_chipselect -> pio_output:chipselect
	signal mm_interconnect_0_pio_output_s1_write                          : std_logic;                     -- mm_interconnect_0:pio_output_s1_write -> mm_interconnect_0_pio_output_s1_write:in
	signal mm_interconnect_0_pio_output_s1_readdata                       : std_logic_vector(31 downto 0); -- pio_output:readdata -> mm_interconnect_0:pio_output_s1_readdata
	signal i2c_master_d_avalon_slave_0_waitrequest                        : std_logic;                     -- i2c_master_d:wb_ack_o -> i2c_master_d_avalon_slave_0_waitrequest:in
	signal mm_interconnect_0_i2c_master_d_avalon_slave_0_writedata        : std_logic_vector(7 downto 0);  -- mm_interconnect_0:i2c_master_d_avalon_slave_0_writedata -> i2c_master_d:wb_dat_i
	signal mm_interconnect_0_i2c_master_d_avalon_slave_0_address          : std_logic_vector(2 downto 0);  -- mm_interconnect_0:i2c_master_d_avalon_slave_0_address -> i2c_master_d:wb_adr_i
	signal mm_interconnect_0_i2c_master_d_avalon_slave_0_chipselect       : std_logic;                     -- mm_interconnect_0:i2c_master_d_avalon_slave_0_chipselect -> i2c_master_d:wb_stb_i
	signal mm_interconnect_0_i2c_master_d_avalon_slave_0_write            : std_logic;                     -- mm_interconnect_0:i2c_master_d_avalon_slave_0_write -> i2c_master_d:wb_we_i
	signal mm_interconnect_0_i2c_master_d_avalon_slave_0_readdata         : std_logic_vector(7 downto 0);  -- i2c_master_d:wb_dat_o -> mm_interconnect_0:i2c_master_d_avalon_slave_0_readdata
	signal i2c_master_f_avalon_slave_0_waitrequest                        : std_logic;                     -- i2c_master_f:wb_ack_o -> i2c_master_f_avalon_slave_0_waitrequest:in
	signal mm_interconnect_0_i2c_master_f_avalon_slave_0_writedata        : std_logic_vector(7 downto 0);  -- mm_interconnect_0:i2c_master_f_avalon_slave_0_writedata -> i2c_master_f:wb_dat_i
	signal mm_interconnect_0_i2c_master_f_avalon_slave_0_address          : std_logic_vector(2 downto 0);  -- mm_interconnect_0:i2c_master_f_avalon_slave_0_address -> i2c_master_f:wb_adr_i
	signal mm_interconnect_0_i2c_master_f_avalon_slave_0_chipselect       : std_logic;                     -- mm_interconnect_0:i2c_master_f_avalon_slave_0_chipselect -> i2c_master_f:wb_stb_i
	signal mm_interconnect_0_i2c_master_f_avalon_slave_0_write            : std_logic;                     -- mm_interconnect_0:i2c_master_f_avalon_slave_0_write -> i2c_master_f:wb_we_i
	signal mm_interconnect_0_i2c_master_f_avalon_slave_0_readdata         : std_logic_vector(7 downto 0);  -- i2c_master_f:wb_dat_o -> mm_interconnect_0:i2c_master_f_avalon_slave_0_readdata
	signal i2c_master_p_avalon_slave_0_waitrequest                        : std_logic;                     -- i2c_master_p:wb_ack_o -> i2c_master_p_avalon_slave_0_waitrequest:in
	signal mm_interconnect_0_i2c_master_p_avalon_slave_0_writedata        : std_logic_vector(7 downto 0);  -- mm_interconnect_0:i2c_master_p_avalon_slave_0_writedata -> i2c_master_p:wb_dat_i
	signal mm_interconnect_0_i2c_master_p_avalon_slave_0_address          : std_logic_vector(2 downto 0);  -- mm_interconnect_0:i2c_master_p_avalon_slave_0_address -> i2c_master_p:wb_adr_i
	signal mm_interconnect_0_i2c_master_p_avalon_slave_0_chipselect       : std_logic;                     -- mm_interconnect_0:i2c_master_p_avalon_slave_0_chipselect -> i2c_master_p:wb_stb_i
	signal mm_interconnect_0_i2c_master_p_avalon_slave_0_write            : std_logic;                     -- mm_interconnect_0:i2c_master_p_avalon_slave_0_write -> i2c_master_p:wb_we_i
	signal mm_interconnect_0_i2c_master_p_avalon_slave_0_readdata         : std_logic_vector(7 downto 0);  -- i2c_master_p:wb_dat_o -> mm_interconnect_0:i2c_master_p_avalon_slave_0_readdata
	signal hps_0_h2f_axi_master_awvalid                                   : std_logic;                     -- hps_0:h2f_AWVALID -> mm_interconnect_1:hps_0_h2f_axi_master_awvalid
	signal hps_0_h2f_axi_master_arsize                                    : std_logic_vector(2 downto 0);  -- hps_0:h2f_ARSIZE -> mm_interconnect_1:hps_0_h2f_axi_master_arsize
	signal hps_0_h2f_axi_master_arlock                                    : std_logic_vector(1 downto 0);  -- hps_0:h2f_ARLOCK -> mm_interconnect_1:hps_0_h2f_axi_master_arlock
	signal hps_0_h2f_axi_master_awcache                                   : std_logic_vector(3 downto 0);  -- hps_0:h2f_AWCACHE -> mm_interconnect_1:hps_0_h2f_axi_master_awcache
	signal hps_0_h2f_axi_master_arready                                   : std_logic;                     -- mm_interconnect_1:hps_0_h2f_axi_master_arready -> hps_0:h2f_ARREADY
	signal hps_0_h2f_axi_master_arid                                      : std_logic_vector(11 downto 0); -- hps_0:h2f_ARID -> mm_interconnect_1:hps_0_h2f_axi_master_arid
	signal hps_0_h2f_axi_master_rready                                    : std_logic;                     -- hps_0:h2f_RREADY -> mm_interconnect_1:hps_0_h2f_axi_master_rready
	signal hps_0_h2f_axi_master_bready                                    : std_logic;                     -- hps_0:h2f_BREADY -> mm_interconnect_1:hps_0_h2f_axi_master_bready
	signal hps_0_h2f_axi_master_awsize                                    : std_logic_vector(2 downto 0);  -- hps_0:h2f_AWSIZE -> mm_interconnect_1:hps_0_h2f_axi_master_awsize
	signal hps_0_h2f_axi_master_awprot                                    : std_logic_vector(2 downto 0);  -- hps_0:h2f_AWPROT -> mm_interconnect_1:hps_0_h2f_axi_master_awprot
	signal hps_0_h2f_axi_master_arvalid                                   : std_logic;                     -- hps_0:h2f_ARVALID -> mm_interconnect_1:hps_0_h2f_axi_master_arvalid
	signal hps_0_h2f_axi_master_arprot                                    : std_logic_vector(2 downto 0);  -- hps_0:h2f_ARPROT -> mm_interconnect_1:hps_0_h2f_axi_master_arprot
	signal hps_0_h2f_axi_master_bid                                       : std_logic_vector(11 downto 0); -- mm_interconnect_1:hps_0_h2f_axi_master_bid -> hps_0:h2f_BID
	signal hps_0_h2f_axi_master_arlen                                     : std_logic_vector(3 downto 0);  -- hps_0:h2f_ARLEN -> mm_interconnect_1:hps_0_h2f_axi_master_arlen
	signal hps_0_h2f_axi_master_awready                                   : std_logic;                     -- mm_interconnect_1:hps_0_h2f_axi_master_awready -> hps_0:h2f_AWREADY
	signal hps_0_h2f_axi_master_awid                                      : std_logic_vector(11 downto 0); -- hps_0:h2f_AWID -> mm_interconnect_1:hps_0_h2f_axi_master_awid
	signal hps_0_h2f_axi_master_bvalid                                    : std_logic;                     -- mm_interconnect_1:hps_0_h2f_axi_master_bvalid -> hps_0:h2f_BVALID
	signal hps_0_h2f_axi_master_wid                                       : std_logic_vector(11 downto 0); -- hps_0:h2f_WID -> mm_interconnect_1:hps_0_h2f_axi_master_wid
	signal hps_0_h2f_axi_master_awlock                                    : std_logic_vector(1 downto 0);  -- hps_0:h2f_AWLOCK -> mm_interconnect_1:hps_0_h2f_axi_master_awlock
	signal hps_0_h2f_axi_master_awburst                                   : std_logic_vector(1 downto 0);  -- hps_0:h2f_AWBURST -> mm_interconnect_1:hps_0_h2f_axi_master_awburst
	signal hps_0_h2f_axi_master_bresp                                     : std_logic_vector(1 downto 0);  -- mm_interconnect_1:hps_0_h2f_axi_master_bresp -> hps_0:h2f_BRESP
	signal hps_0_h2f_axi_master_wstrb                                     : std_logic_vector(7 downto 0);  -- hps_0:h2f_WSTRB -> mm_interconnect_1:hps_0_h2f_axi_master_wstrb
	signal hps_0_h2f_axi_master_rvalid                                    : std_logic;                     -- mm_interconnect_1:hps_0_h2f_axi_master_rvalid -> hps_0:h2f_RVALID
	signal hps_0_h2f_axi_master_wdata                                     : std_logic_vector(63 downto 0); -- hps_0:h2f_WDATA -> mm_interconnect_1:hps_0_h2f_axi_master_wdata
	signal hps_0_h2f_axi_master_wready                                    : std_logic;                     -- mm_interconnect_1:hps_0_h2f_axi_master_wready -> hps_0:h2f_WREADY
	signal hps_0_h2f_axi_master_arburst                                   : std_logic_vector(1 downto 0);  -- hps_0:h2f_ARBURST -> mm_interconnect_1:hps_0_h2f_axi_master_arburst
	signal hps_0_h2f_axi_master_rdata                                     : std_logic_vector(63 downto 0); -- mm_interconnect_1:hps_0_h2f_axi_master_rdata -> hps_0:h2f_RDATA
	signal hps_0_h2f_axi_master_araddr                                    : std_logic_vector(29 downto 0); -- hps_0:h2f_ARADDR -> mm_interconnect_1:hps_0_h2f_axi_master_araddr
	signal hps_0_h2f_axi_master_arcache                                   : std_logic_vector(3 downto 0);  -- hps_0:h2f_ARCACHE -> mm_interconnect_1:hps_0_h2f_axi_master_arcache
	signal hps_0_h2f_axi_master_awlen                                     : std_logic_vector(3 downto 0);  -- hps_0:h2f_AWLEN -> mm_interconnect_1:hps_0_h2f_axi_master_awlen
	signal hps_0_h2f_axi_master_awaddr                                    : std_logic_vector(29 downto 0); -- hps_0:h2f_AWADDR -> mm_interconnect_1:hps_0_h2f_axi_master_awaddr
	signal hps_0_h2f_axi_master_rid                                       : std_logic_vector(11 downto 0); -- mm_interconnect_1:hps_0_h2f_axi_master_rid -> hps_0:h2f_RID
	signal hps_0_h2f_axi_master_wvalid                                    : std_logic;                     -- hps_0:h2f_WVALID -> mm_interconnect_1:hps_0_h2f_axi_master_wvalid
	signal hps_0_h2f_axi_master_rresp                                     : std_logic_vector(1 downto 0);  -- mm_interconnect_1:hps_0_h2f_axi_master_rresp -> hps_0:h2f_RRESP
	signal hps_0_h2f_axi_master_wlast                                     : std_logic;                     -- hps_0:h2f_WLAST -> mm_interconnect_1:hps_0_h2f_axi_master_wlast
	signal hps_0_h2f_axi_master_rlast                                     : std_logic;                     -- mm_interconnect_1:hps_0_h2f_axi_master_rlast -> hps_0:h2f_RLAST
	signal mm_interconnect_1_sld_hub_controller_system_0_s0_waitrequest   : std_logic;                     -- sld_hub_controller_system_0:s0_waitrequest -> mm_interconnect_1:sld_hub_controller_system_0_s0_waitrequest
	signal mm_interconnect_1_sld_hub_controller_system_0_s0_burstcount    : std_logic_vector(0 downto 0);  -- mm_interconnect_1:sld_hub_controller_system_0_s0_burstcount -> sld_hub_controller_system_0:s0_burstcount
	signal mm_interconnect_1_sld_hub_controller_system_0_s0_writedata     : std_logic_vector(31 downto 0); -- mm_interconnect_1:sld_hub_controller_system_0_s0_writedata -> sld_hub_controller_system_0:s0_writedata
	signal mm_interconnect_1_sld_hub_controller_system_0_s0_address       : std_logic_vector(6 downto 0);  -- mm_interconnect_1:sld_hub_controller_system_0_s0_address -> sld_hub_controller_system_0:s0_address
	signal mm_interconnect_1_sld_hub_controller_system_0_s0_write         : std_logic;                     -- mm_interconnect_1:sld_hub_controller_system_0_s0_write -> sld_hub_controller_system_0:s0_write
	signal mm_interconnect_1_sld_hub_controller_system_0_s0_read          : std_logic;                     -- mm_interconnect_1:sld_hub_controller_system_0_s0_read -> sld_hub_controller_system_0:s0_read
	signal mm_interconnect_1_sld_hub_controller_system_0_s0_readdata      : std_logic_vector(31 downto 0); -- sld_hub_controller_system_0:s0_readdata -> mm_interconnect_1:sld_hub_controller_system_0_s0_readdata
	signal mm_interconnect_1_sld_hub_controller_system_0_s0_debugaccess   : std_logic;                     -- mm_interconnect_1:sld_hub_controller_system_0_s0_debugaccess -> sld_hub_controller_system_0:s0_debugaccess
	signal mm_interconnect_1_sld_hub_controller_system_0_s0_readdatavalid : std_logic;                     -- sld_hub_controller_system_0:s0_readdatavalid -> mm_interconnect_1:sld_hub_controller_system_0_s0_readdatavalid
	signal mm_interconnect_1_sld_hub_controller_system_0_s0_byteenable    : std_logic_vector(3 downto 0);  -- mm_interconnect_1:sld_hub_controller_system_0_s0_byteenable -> sld_hub_controller_system_0:s0_byteenable
	signal mm_interconnect_1_onchip_memory_nios_cpu_s2_writedata          : std_logic_vector(31 downto 0); -- mm_interconnect_1:onchip_memory_nios_cpu_s2_writedata -> onchip_memory_nios_cpu:writedata2
	signal mm_interconnect_1_onchip_memory_nios_cpu_s2_address            : std_logic_vector(13 downto 0); -- mm_interconnect_1:onchip_memory_nios_cpu_s2_address -> onchip_memory_nios_cpu:address2
	signal mm_interconnect_1_onchip_memory_nios_cpu_s2_chipselect         : std_logic;                     -- mm_interconnect_1:onchip_memory_nios_cpu_s2_chipselect -> onchip_memory_nios_cpu:chipselect2
	signal mm_interconnect_1_onchip_memory_nios_cpu_s2_clken              : std_logic;                     -- mm_interconnect_1:onchip_memory_nios_cpu_s2_clken -> onchip_memory_nios_cpu:clken2
	signal mm_interconnect_1_onchip_memory_nios_cpu_s2_write              : std_logic;                     -- mm_interconnect_1:onchip_memory_nios_cpu_s2_write -> onchip_memory_nios_cpu:write2
	signal mm_interconnect_1_onchip_memory_nios_cpu_s2_readdata           : std_logic_vector(31 downto 0); -- onchip_memory_nios_cpu:readdata2 -> mm_interconnect_1:onchip_memory_nios_cpu_s2_readdata
	signal mm_interconnect_1_onchip_memory_nios_cpu_s2_byteenable         : std_logic_vector(3 downto 0);  -- mm_interconnect_1:onchip_memory_nios_cpu_s2_byteenable -> onchip_memory_nios_cpu:byteenable2
	signal mm_interconnect_1_onchip_memory_nios_arm_s2_writedata          : std_logic_vector(15 downto 0); -- mm_interconnect_1:onchip_memory_nios_arm_s2_writedata -> onchip_memory_nios_arm:writedata2
	signal mm_interconnect_1_onchip_memory_nios_arm_s2_address            : std_logic_vector(14 downto 0); -- mm_interconnect_1:onchip_memory_nios_arm_s2_address -> onchip_memory_nios_arm:address2
	signal mm_interconnect_1_onchip_memory_nios_arm_s2_chipselect         : std_logic;                     -- mm_interconnect_1:onchip_memory_nios_arm_s2_chipselect -> onchip_memory_nios_arm:chipselect2
	signal mm_interconnect_1_onchip_memory_nios_arm_s2_clken              : std_logic;                     -- mm_interconnect_1:onchip_memory_nios_arm_s2_clken -> onchip_memory_nios_arm:clken2
	signal mm_interconnect_1_onchip_memory_nios_arm_s2_write              : std_logic;                     -- mm_interconnect_1:onchip_memory_nios_arm_s2_write -> onchip_memory_nios_arm:write2
	signal mm_interconnect_1_onchip_memory_nios_arm_s2_readdata           : std_logic_vector(15 downto 0); -- onchip_memory_nios_arm:readdata2 -> mm_interconnect_1:onchip_memory_nios_arm_s2_readdata
	signal mm_interconnect_1_onchip_memory_nios_arm_s2_byteenable         : std_logic_vector(1 downto 0);  -- mm_interconnect_1:onchip_memory_nios_arm_s2_byteenable -> onchip_memory_nios_arm:byteenable2
	signal hps_0_f2h_irq0_irq                                             : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> hps_0:f2h_irq_p0
	signal hps_0_f2h_irq1_irq                                             : std_logic_vector(31 downto 0); -- irq_mapper_001:sender_irq -> hps_0:f2h_irq_p1
	signal irq_mapper_002_receiver0_irq                                   : std_logic;                     -- timer_0:irq -> irq_mapper_002:receiver0_irq
	signal irq_mapper_002_receiver1_irq                                   : std_logic;                     -- timer_1:irq -> irq_mapper_002:receiver1_irq
	signal irq_mapper_002_receiver2_irq                                   : std_logic;                     -- i2c_master_is1:wb_inta_o -> irq_mapper_002:receiver2_irq
	signal irq_mapper_002_receiver3_irq                                   : std_logic;                     -- i2c_master_is2:wb_inta_o -> irq_mapper_002:receiver3_irq
	signal irq_mapper_002_receiver4_irq                                   : std_logic;                     -- i2c_master_is3:wb_inta_o -> irq_mapper_002:receiver4_irq
	signal irq_mapper_002_receiver5_irq                                   : std_logic;                     -- i2c_master_is4:wb_inta_o -> irq_mapper_002:receiver5_irq
	signal irq_mapper_002_receiver6_irq                                   : std_logic;                     -- pio_input:irq -> irq_mapper_002:receiver6_irq
	signal irq_mapper_002_receiver8_irq                                   : std_logic;                     -- i2c_master_d:wb_inta_o -> irq_mapper_002:receiver8_irq
	signal irq_mapper_002_receiver9_irq                                   : std_logic;                     -- i2c_master_f:wb_inta_o -> irq_mapper_002:receiver9_irq
	signal irq_mapper_002_receiver10_irq                                  : std_logic;                     -- i2c_master_p:wb_inta_o -> irq_mapper_002:receiver10_irq
	signal nios2_qsys_0_d_irq_irq                                         : std_logic_vector(31 downto 0); -- irq_mapper_002:sender_irq -> nios2_qsys_0:d_irq
	signal irq_mapper_receiver0_irq                                       : std_logic;                     -- jtag_uart:av_irq -> [irq_mapper:receiver0_irq, irq_mapper_002:receiver7_irq]
	signal rst_controller_reset_out_reset                                 : std_logic;                     -- rst_controller:reset_out -> [mm_interconnect_0:sysid_reset_reset_bridge_in_reset_reset, mm_interconnect_1:sld_hub_controller_system_0_reset_reset_bridge_in_reset_reset, onchip_memory_nios_arm:reset, onchip_memory_nios_cpu:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset, sld_hub_controller_system_0:reset_reset]
	signal rst_controller_reset_out_reset_req                             : std_logic;                     -- rst_controller:reset_req -> [onchip_memory_nios_arm:reset_req, onchip_memory_nios_cpu:reset_req, rst_translator:reset_req_in]
	signal hps_0_h2f_reset_reset                                          : std_logic;                     -- hps_0:h2f_rst_n -> hps_0_h2f_reset_reset:in
	signal rst_controller_001_reset_out_reset                             : std_logic;                     -- rst_controller_001:reset_out -> [i2c_master_d:wb_rst_i, i2c_master_f:wb_rst_i, i2c_master_is1:wb_rst_i, i2c_master_is2:wb_rst_i, i2c_master_is3:wb_rst_i, i2c_master_is4:wb_rst_i, i2c_master_p:wb_rst_i, irq_mapper_002:reset, mm_interconnect_0:fpga_only_master_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_0:nios2_qsys_0_reset_n_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in, rst_translator_001:in_reset]
	signal rst_controller_001_reset_out_reset_req                         : std_logic;                     -- rst_controller_001:reset_req -> [nios2_qsys_0:reset_req, rst_translator_001:reset_req_in]
	signal rst_controller_002_reset_out_reset                             : std_logic;                     -- rst_controller_002:reset_out -> [mm_interconnect_0:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset]
	signal qsys_reset_reset_n_ports_inv                                   : std_logic;                     -- qsys_reset_reset_n:inv -> [fpga_only_master:clk_reset_reset, rst_controller:reset_in1, rst_controller_001:reset_in0]
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv   : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_0_pio_reset_nios_s1_write_ports_inv            : std_logic;                     -- mm_interconnect_0_pio_reset_nios_s1_write:inv -> pio_reset_nios:write_n
	signal mm_interconnect_0_timer_0_s1_write_ports_inv                   : std_logic;                     -- mm_interconnect_0_timer_0_s1_write:inv -> timer_0:write_n
	signal mm_interconnect_0_timer_1_s1_write_ports_inv                   : std_logic;                     -- mm_interconnect_0_timer_1_s1_write:inv -> timer_1:write_n
	signal mm_interconnect_0_i2c_master_is1_avalon_slave_0_inv            : std_logic;                     -- i2c_master_is1_avalon_slave_0_waitrequest:inv -> mm_interconnect_0:i2c_master_is1_avalon_slave_0_waitrequest
	signal mm_interconnect_0_i2c_master_is2_avalon_slave_0_inv            : std_logic;                     -- i2c_master_is2_avalon_slave_0_waitrequest:inv -> mm_interconnect_0:i2c_master_is2_avalon_slave_0_waitrequest
	signal mm_interconnect_0_i2c_master_is3_avalon_slave_0_inv            : std_logic;                     -- i2c_master_is3_avalon_slave_0_waitrequest:inv -> mm_interconnect_0:i2c_master_is3_avalon_slave_0_waitrequest
	signal mm_interconnect_0_i2c_master_is4_avalon_slave_0_inv            : std_logic;                     -- i2c_master_is4_avalon_slave_0_waitrequest:inv -> mm_interconnect_0:i2c_master_is4_avalon_slave_0_waitrequest
	signal mm_interconnect_0_pio_input_s1_write_ports_inv                 : std_logic;                     -- mm_interconnect_0_pio_input_s1_write:inv -> pio_input:write_n
	signal mm_interconnect_0_pio_output_s1_write_ports_inv                : std_logic;                     -- mm_interconnect_0_pio_output_s1_write:inv -> pio_output:write_n
	signal mm_interconnect_0_i2c_master_d_avalon_slave_0_inv              : std_logic;                     -- i2c_master_d_avalon_slave_0_waitrequest:inv -> mm_interconnect_0:i2c_master_d_avalon_slave_0_waitrequest
	signal mm_interconnect_0_i2c_master_f_avalon_slave_0_inv              : std_logic;                     -- i2c_master_f_avalon_slave_0_waitrequest:inv -> mm_interconnect_0:i2c_master_f_avalon_slave_0_waitrequest
	signal mm_interconnect_0_i2c_master_p_avalon_slave_0_inv              : std_logic;                     -- i2c_master_p_avalon_slave_0_waitrequest:inv -> mm_interconnect_0:i2c_master_p_avalon_slave_0_waitrequest
	signal rst_controller_reset_out_reset_ports_inv                       : std_logic;                     -- rst_controller_reset_out_reset:inv -> [pio_reset_nios:reset_n, sysid:reset_n]
	signal hps_0_h2f_reset_reset_ports_inv                                : std_logic;                     -- hps_0_h2f_reset_reset:inv -> [rst_controller:reset_in0, rst_controller_002:reset_in0]
	signal rst_controller_001_reset_out_reset_ports_inv                   : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> [avalon_spi_AMC7891_0:csi_clock_reset_n, avalon_spi_AMC7891_1:csi_clock_reset_n, jtag_uart:rst_n, nios2_qsys_0:reset_n, pio_input:reset_n, pio_output:reset_n, timer_0:reset_n, timer_1:reset_n]

begin

	hps_0 : component fluid_board_soc_hps_0
		generic map (
			F2S_Width => 0,
			S2F_Width => 2
		)
		port map (
			uart1_cts                => hps_0_uart1_cts,                 --             uart1.cts
			uart1_dsr                => hps_0_uart1_dsr,                 --                  .dsr
			uart1_dcd                => hps_0_uart1_dcd,                 --                  .dcd
			uart1_ri                 => hps_0_uart1_ri,                  --                  .ri
			uart1_dtr                => hps_0_uart1_dtr,                 --                  .dtr
			uart1_rts                => hps_0_uart1_rts,                 --                  .rts
			uart1_out1_n             => hps_0_uart1_out1_n,              --                  .out1_n
			uart1_out2_n             => hps_0_uart1_out2_n,              --                  .out2_n
			uart1_rxd                => hps_0_uart1_rxd,                 --                  .rxd
			uart1_txd                => hps_0_uart1_txd,                 --                  .txd
			mem_a                    => memory_mem_a,                    --            memory.mem_a
			mem_ba                   => memory_mem_ba,                   --                  .mem_ba
			mem_ck                   => memory_mem_ck,                   --                  .mem_ck
			mem_ck_n                 => memory_mem_ck_n,                 --                  .mem_ck_n
			mem_cke                  => memory_mem_cke,                  --                  .mem_cke
			mem_cs_n                 => memory_mem_cs_n,                 --                  .mem_cs_n
			mem_ras_n                => memory_mem_ras_n,                --                  .mem_ras_n
			mem_cas_n                => memory_mem_cas_n,                --                  .mem_cas_n
			mem_we_n                 => memory_mem_we_n,                 --                  .mem_we_n
			mem_reset_n              => memory_mem_reset_n,              --                  .mem_reset_n
			mem_dq                   => memory_mem_dq,                   --                  .mem_dq
			mem_dqs                  => memory_mem_dqs,                  --                  .mem_dqs
			mem_dqs_n                => memory_mem_dqs_n,                --                  .mem_dqs_n
			mem_odt                  => memory_mem_odt,                  --                  .mem_odt
			mem_dm                   => memory_mem_dm,                   --                  .mem_dm
			oct_rzqin                => memory_oct_rzqin,                --                  .oct_rzqin
			hps_io_emac0_inst_TX_CLK => hps_io_hps_io_emac0_inst_TX_CLK, --            hps_io.hps_io_emac0_inst_TX_CLK
			hps_io_emac0_inst_TXD0   => hps_io_hps_io_emac0_inst_TXD0,   --                  .hps_io_emac0_inst_TXD0
			hps_io_emac0_inst_TXD1   => hps_io_hps_io_emac0_inst_TXD1,   --                  .hps_io_emac0_inst_TXD1
			hps_io_emac0_inst_TXD2   => hps_io_hps_io_emac0_inst_TXD2,   --                  .hps_io_emac0_inst_TXD2
			hps_io_emac0_inst_TXD3   => hps_io_hps_io_emac0_inst_TXD3,   --                  .hps_io_emac0_inst_TXD3
			hps_io_emac0_inst_RXD0   => hps_io_hps_io_emac0_inst_RXD0,   --                  .hps_io_emac0_inst_RXD0
			hps_io_emac0_inst_MDIO   => hps_io_hps_io_emac0_inst_MDIO,   --                  .hps_io_emac0_inst_MDIO
			hps_io_emac0_inst_MDC    => hps_io_hps_io_emac0_inst_MDC,    --                  .hps_io_emac0_inst_MDC
			hps_io_emac0_inst_RX_CTL => hps_io_hps_io_emac0_inst_RX_CTL, --                  .hps_io_emac0_inst_RX_CTL
			hps_io_emac0_inst_TX_CTL => hps_io_hps_io_emac0_inst_TX_CTL, --                  .hps_io_emac0_inst_TX_CTL
			hps_io_emac0_inst_RX_CLK => hps_io_hps_io_emac0_inst_RX_CLK, --                  .hps_io_emac0_inst_RX_CLK
			hps_io_emac0_inst_RXD1   => hps_io_hps_io_emac0_inst_RXD1,   --                  .hps_io_emac0_inst_RXD1
			hps_io_emac0_inst_RXD2   => hps_io_hps_io_emac0_inst_RXD2,   --                  .hps_io_emac0_inst_RXD2
			hps_io_emac0_inst_RXD3   => hps_io_hps_io_emac0_inst_RXD3,   --                  .hps_io_emac0_inst_RXD3
			hps_io_uart0_inst_RX     => hps_io_hps_io_uart0_inst_RX,     --                  .hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX     => hps_io_hps_io_uart0_inst_TX,     --                  .hps_io_uart0_inst_TX
			hps_io_gpio_inst_GPIO26  => hps_io_hps_io_gpio_inst_GPIO26,  --                  .hps_io_gpio_inst_GPIO26
			hps_io_gpio_inst_GPIO28  => hps_io_hps_io_gpio_inst_GPIO28,  --                  .hps_io_gpio_inst_GPIO28
			hps_io_gpio_inst_GPIO59  => hps_io_hps_io_gpio_inst_GPIO59,  --                  .hps_io_gpio_inst_GPIO59
			h2f_rst_n                => hps_0_h2f_reset_reset,           --         h2f_reset.reset_n
			h2f_axi_clk              => pll_0_outclk0_clk,               --     h2f_axi_clock.clk
			h2f_AWID                 => hps_0_h2f_axi_master_awid,       --    h2f_axi_master.awid
			h2f_AWADDR               => hps_0_h2f_axi_master_awaddr,     --                  .awaddr
			h2f_AWLEN                => hps_0_h2f_axi_master_awlen,      --                  .awlen
			h2f_AWSIZE               => hps_0_h2f_axi_master_awsize,     --                  .awsize
			h2f_AWBURST              => hps_0_h2f_axi_master_awburst,    --                  .awburst
			h2f_AWLOCK               => hps_0_h2f_axi_master_awlock,     --                  .awlock
			h2f_AWCACHE              => hps_0_h2f_axi_master_awcache,    --                  .awcache
			h2f_AWPROT               => hps_0_h2f_axi_master_awprot,     --                  .awprot
			h2f_AWVALID              => hps_0_h2f_axi_master_awvalid,    --                  .awvalid
			h2f_AWREADY              => hps_0_h2f_axi_master_awready,    --                  .awready
			h2f_WID                  => hps_0_h2f_axi_master_wid,        --                  .wid
			h2f_WDATA                => hps_0_h2f_axi_master_wdata,      --                  .wdata
			h2f_WSTRB                => hps_0_h2f_axi_master_wstrb,      --                  .wstrb
			h2f_WLAST                => hps_0_h2f_axi_master_wlast,      --                  .wlast
			h2f_WVALID               => hps_0_h2f_axi_master_wvalid,     --                  .wvalid
			h2f_WREADY               => hps_0_h2f_axi_master_wready,     --                  .wready
			h2f_BID                  => hps_0_h2f_axi_master_bid,        --                  .bid
			h2f_BRESP                => hps_0_h2f_axi_master_bresp,      --                  .bresp
			h2f_BVALID               => hps_0_h2f_axi_master_bvalid,     --                  .bvalid
			h2f_BREADY               => hps_0_h2f_axi_master_bready,     --                  .bready
			h2f_ARID                 => hps_0_h2f_axi_master_arid,       --                  .arid
			h2f_ARADDR               => hps_0_h2f_axi_master_araddr,     --                  .araddr
			h2f_ARLEN                => hps_0_h2f_axi_master_arlen,      --                  .arlen
			h2f_ARSIZE               => hps_0_h2f_axi_master_arsize,     --                  .arsize
			h2f_ARBURST              => hps_0_h2f_axi_master_arburst,    --                  .arburst
			h2f_ARLOCK               => hps_0_h2f_axi_master_arlock,     --                  .arlock
			h2f_ARCACHE              => hps_0_h2f_axi_master_arcache,    --                  .arcache
			h2f_ARPROT               => hps_0_h2f_axi_master_arprot,     --                  .arprot
			h2f_ARVALID              => hps_0_h2f_axi_master_arvalid,    --                  .arvalid
			h2f_ARREADY              => hps_0_h2f_axi_master_arready,    --                  .arready
			h2f_RID                  => hps_0_h2f_axi_master_rid,        --                  .rid
			h2f_RDATA                => hps_0_h2f_axi_master_rdata,      --                  .rdata
			h2f_RRESP                => hps_0_h2f_axi_master_rresp,      --                  .rresp
			h2f_RLAST                => hps_0_h2f_axi_master_rlast,      --                  .rlast
			h2f_RVALID               => hps_0_h2f_axi_master_rvalid,     --                  .rvalid
			h2f_RREADY               => hps_0_h2f_axi_master_rready,     --                  .rready
			h2f_lw_axi_clk           => pll_0_outclk0_clk,               --  h2f_lw_axi_clock.clk
			h2f_lw_AWID              => hps_0_h2f_lw_axi_master_awid,    -- h2f_lw_axi_master.awid
			h2f_lw_AWADDR            => hps_0_h2f_lw_axi_master_awaddr,  --                  .awaddr
			h2f_lw_AWLEN             => hps_0_h2f_lw_axi_master_awlen,   --                  .awlen
			h2f_lw_AWSIZE            => hps_0_h2f_lw_axi_master_awsize,  --                  .awsize
			h2f_lw_AWBURST           => hps_0_h2f_lw_axi_master_awburst, --                  .awburst
			h2f_lw_AWLOCK            => hps_0_h2f_lw_axi_master_awlock,  --                  .awlock
			h2f_lw_AWCACHE           => hps_0_h2f_lw_axi_master_awcache, --                  .awcache
			h2f_lw_AWPROT            => hps_0_h2f_lw_axi_master_awprot,  --                  .awprot
			h2f_lw_AWVALID           => hps_0_h2f_lw_axi_master_awvalid, --                  .awvalid
			h2f_lw_AWREADY           => hps_0_h2f_lw_axi_master_awready, --                  .awready
			h2f_lw_WID               => hps_0_h2f_lw_axi_master_wid,     --                  .wid
			h2f_lw_WDATA             => hps_0_h2f_lw_axi_master_wdata,   --                  .wdata
			h2f_lw_WSTRB             => hps_0_h2f_lw_axi_master_wstrb,   --                  .wstrb
			h2f_lw_WLAST             => hps_0_h2f_lw_axi_master_wlast,   --                  .wlast
			h2f_lw_WVALID            => hps_0_h2f_lw_axi_master_wvalid,  --                  .wvalid
			h2f_lw_WREADY            => hps_0_h2f_lw_axi_master_wready,  --                  .wready
			h2f_lw_BID               => hps_0_h2f_lw_axi_master_bid,     --                  .bid
			h2f_lw_BRESP             => hps_0_h2f_lw_axi_master_bresp,   --                  .bresp
			h2f_lw_BVALID            => hps_0_h2f_lw_axi_master_bvalid,  --                  .bvalid
			h2f_lw_BREADY            => hps_0_h2f_lw_axi_master_bready,  --                  .bready
			h2f_lw_ARID              => hps_0_h2f_lw_axi_master_arid,    --                  .arid
			h2f_lw_ARADDR            => hps_0_h2f_lw_axi_master_araddr,  --                  .araddr
			h2f_lw_ARLEN             => hps_0_h2f_lw_axi_master_arlen,   --                  .arlen
			h2f_lw_ARSIZE            => hps_0_h2f_lw_axi_master_arsize,  --                  .arsize
			h2f_lw_ARBURST           => hps_0_h2f_lw_axi_master_arburst, --                  .arburst
			h2f_lw_ARLOCK            => hps_0_h2f_lw_axi_master_arlock,  --                  .arlock
			h2f_lw_ARCACHE           => hps_0_h2f_lw_axi_master_arcache, --                  .arcache
			h2f_lw_ARPROT            => hps_0_h2f_lw_axi_master_arprot,  --                  .arprot
			h2f_lw_ARVALID           => hps_0_h2f_lw_axi_master_arvalid, --                  .arvalid
			h2f_lw_ARREADY           => hps_0_h2f_lw_axi_master_arready, --                  .arready
			h2f_lw_RID               => hps_0_h2f_lw_axi_master_rid,     --                  .rid
			h2f_lw_RDATA             => hps_0_h2f_lw_axi_master_rdata,   --                  .rdata
			h2f_lw_RRESP             => hps_0_h2f_lw_axi_master_rresp,   --                  .rresp
			h2f_lw_RLAST             => hps_0_h2f_lw_axi_master_rlast,   --                  .rlast
			h2f_lw_RVALID            => hps_0_h2f_lw_axi_master_rvalid,  --                  .rvalid
			h2f_lw_RREADY            => hps_0_h2f_lw_axi_master_rready,  --                  .rready
			f2h_irq_p0               => hps_0_f2h_irq0_irq,              --          f2h_irq0.irq
			f2h_irq_p1               => hps_0_f2h_irq1_irq               --          f2h_irq1.irq
		);

	sysid : component fluid_board_soc_sysid
		port map (
			clock    => pll_0_outclk0_clk,                                --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,         --         reset.reset_n
			readdata => mm_interconnect_0_sysid_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_control_slave_address(0)  --              .address
		);

	pll_0 : component fluid_board_soc_pll_0
		port map (
			refclk   => pll_0_refclk_clk,    --  refclk.clk
			rst      => pll_0_reset_reset,   --   reset.reset
			outclk_0 => pll_0_outclk0_clk,   -- outclk0.clk
			locked   => pll_0_locked_export  --  locked.export
		);

	sld_hub_controller_system_0 : component fluid_board_soc_sld_hub_controller_system_0
		generic map (
			ENABLE_JTAG_IO_SELECTION => 0
		)
		port map (
			clk_clk          => pll_0_outclk0_clk,                                              --   clk.clk
			reset_reset      => rst_controller_reset_out_reset,                                 -- reset.reset
			s0_waitrequest   => mm_interconnect_1_sld_hub_controller_system_0_s0_waitrequest,   --    s0.waitrequest
			s0_readdata      => mm_interconnect_1_sld_hub_controller_system_0_s0_readdata,      --      .readdata
			s0_readdatavalid => mm_interconnect_1_sld_hub_controller_system_0_s0_readdatavalid, --      .readdatavalid
			s0_burstcount    => mm_interconnect_1_sld_hub_controller_system_0_s0_burstcount,    --      .burstcount
			s0_writedata     => mm_interconnect_1_sld_hub_controller_system_0_s0_writedata,     --      .writedata
			s0_address       => mm_interconnect_1_sld_hub_controller_system_0_s0_address,       --      .address
			s0_write         => mm_interconnect_1_sld_hub_controller_system_0_s0_write,         --      .write
			s0_read          => mm_interconnect_1_sld_hub_controller_system_0_s0_read,          --      .read
			s0_byteenable    => mm_interconnect_1_sld_hub_controller_system_0_s0_byteenable,    --      .byteenable
			s0_debugaccess   => mm_interconnect_1_sld_hub_controller_system_0_s0_debugaccess    --      .debugaccess
		);

	nios2_qsys_0 : component fluid_board_soc_nios2_qsys_0
		port map (
			clk                                   => pll_0_outclk0_clk,                                            --                       clk.clk
			reset_n                               => rst_controller_001_reset_out_reset_ports_inv,                 --                   reset_n.reset_n
			reset_req                             => rst_controller_001_reset_out_reset_req,                       --                          .reset_req
			d_address                             => nios2_qsys_0_data_master_address,                             --               data_master.address
			d_byteenable                          => nios2_qsys_0_data_master_byteenable,                          --                          .byteenable
			d_read                                => nios2_qsys_0_data_master_read,                                --                          .read
			d_readdata                            => nios2_qsys_0_data_master_readdata,                            --                          .readdata
			d_waitrequest                         => nios2_qsys_0_data_master_waitrequest,                         --                          .waitrequest
			d_write                               => nios2_qsys_0_data_master_write,                               --                          .write
			d_writedata                           => nios2_qsys_0_data_master_writedata,                           --                          .writedata
			jtag_debug_module_debugaccess_to_roms => nios2_qsys_0_data_master_debugaccess,                         --                          .debugaccess
			i_address                             => nios2_qsys_0_instruction_master_address,                      --        instruction_master.address
			i_read                                => nios2_qsys_0_instruction_master_read,                         --                          .read
			i_readdata                            => nios2_qsys_0_instruction_master_readdata,                     --                          .readdata
			i_waitrequest                         => nios2_qsys_0_instruction_master_waitrequest,                  --                          .waitrequest
			i_readdatavalid                       => nios2_qsys_0_instruction_master_readdatavalid,                --                          .readdatavalid
			d_irq                                 => nios2_qsys_0_d_irq_irq,                                       --                     d_irq.irq
			jtag_debug_module_resetrequest        => open,                                                         --   jtag_debug_module_reset.reset
			jtag_debug_module_address             => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address,     --         jtag_debug_module.address
			jtag_debug_module_byteenable          => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable,  --                          .byteenable
			jtag_debug_module_debugaccess         => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess, --                          .debugaccess
			jtag_debug_module_read                => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read,        --                          .read
			jtag_debug_module_readdata            => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata,    --                          .readdata
			jtag_debug_module_waitrequest         => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest, --                          .waitrequest
			jtag_debug_module_write               => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write,       --                          .write
			jtag_debug_module_writedata           => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata,   --                          .writedata
			no_ci_readra                          => open,                                                         -- custom_instruction_master.readra
			cpu_resetrequest                      => nios2_qsys_0_cpu_resetrequest_conduit_resetrequest,           --  cpu_resetrequest_conduit.export
			cpu_resettaken                        => nios2_qsys_0_cpu_resetrequest_conduit_resettaken              --                          .export
		);

	timer_0 : component fluid_board_soc_timer_0
		port map (
			clk        => pll_0_outclk0_clk,                            --   clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, -- reset.reset_n
			address    => mm_interconnect_0_timer_0_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_0_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_0_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_0_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_0_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_002_receiver0_irq                  --   irq.irq
		);

	timer_1 : component fluid_board_soc_timer_0
		port map (
			clk        => pll_0_outclk0_clk,                            --   clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, -- reset.reset_n
			address    => mm_interconnect_0_timer_1_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_1_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_1_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_1_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_1_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_002_receiver1_irq                  --   irq.irq
		);

	avalon_spi_amc7891_0 : component avalon_spi_AMC7891
		port map (
			csi_clock_clk      => pll_0_outclk0_clk,                                     --       clock.clk
			csi_clock_reset_n  => rst_controller_001_reset_out_reset_ports_inv,          -- clock_reset.reset_n
			avs_s1_writedata   => mm_interconnect_0_avalon_spi_amc7891_0_s1_writedata,   --          s1.writedata
			avs_s1_read        => mm_interconnect_0_avalon_spi_amc7891_0_s1_read,        --            .read
			avs_s1_write       => mm_interconnect_0_avalon_spi_amc7891_0_s1_write,       --            .write
			avs_s1_address     => mm_interconnect_0_avalon_spi_amc7891_0_s1_address,     --            .address
			avs_s1_waitrequest => mm_interconnect_0_avalon_spi_amc7891_0_s1_waitrequest, --            .waitrequest
			avs_s1_readdata    => mm_interconnect_0_avalon_spi_amc7891_0_s1_readdata,    --            .readdata
			coe_s1_sclk        => avalon_spi_amc7891_0_conduit_end_sclk,                 -- conduit_end.sclk
			coe_s1_cs_n        => avalon_spi_amc7891_0_conduit_end_cs_n,                 --            .cs_n
			coe_s1_sdio        => avalon_spi_amc7891_0_conduit_end_sdio,                 --            .sdio
			coe_s1_sdo         => avalon_spi_amc7891_0_conduit_end_sdo                   --            .sdo
		);

	avalon_spi_amc7891_1 : component avalon_spi_AMC7891
		port map (
			csi_clock_clk      => pll_0_outclk0_clk,                                     --       clock.clk
			csi_clock_reset_n  => rst_controller_001_reset_out_reset_ports_inv,          -- clock_reset.reset_n
			avs_s1_writedata   => mm_interconnect_0_avalon_spi_amc7891_1_s1_writedata,   --          s1.writedata
			avs_s1_read        => mm_interconnect_0_avalon_spi_amc7891_1_s1_read,        --            .read
			avs_s1_write       => mm_interconnect_0_avalon_spi_amc7891_1_s1_write,       --            .write
			avs_s1_address     => mm_interconnect_0_avalon_spi_amc7891_1_s1_address,     --            .address
			avs_s1_waitrequest => mm_interconnect_0_avalon_spi_amc7891_1_s1_waitrequest, --            .waitrequest
			avs_s1_readdata    => mm_interconnect_0_avalon_spi_amc7891_1_s1_readdata,    --            .readdata
			coe_s1_sclk        => avalon_spi_amc7891_1_conduit_end_sclk,                 -- conduit_end.sclk
			coe_s1_cs_n        => avalon_spi_amc7891_1_conduit_end_cs_n,                 --            .cs_n
			coe_s1_sdio        => avalon_spi_amc7891_1_conduit_end_sdio,                 --            .sdio
			coe_s1_sdo         => avalon_spi_amc7891_1_conduit_end_sdo                   --            .sdo
		);

	i2c_master_is1 : component i2c_opencores
		port map (
			wb_adr_i   => mm_interconnect_0_i2c_master_is1_avalon_slave_0_address,    --   avalon_slave_0.address
			wb_dat_i   => mm_interconnect_0_i2c_master_is1_avalon_slave_0_writedata,  --                 .writedata
			wb_dat_o   => mm_interconnect_0_i2c_master_is1_avalon_slave_0_readdata,   --                 .readdata
			wb_we_i    => mm_interconnect_0_i2c_master_is1_avalon_slave_0_write,      --                 .write
			wb_stb_i   => mm_interconnect_0_i2c_master_is1_avalon_slave_0_chipselect, --                 .chipselect
			wb_ack_o   => i2c_master_is1_avalon_slave_0_waitrequest,                  --                 .waitrequest_n
			scl_pad_io => i2c_master_is1_conduit_end_scl,                             --      conduit_end.scl
			sda_pad_io => i2c_master_is1_conduit_end_sda,                             --                 .sda
			wb_clk_i   => pll_0_outclk0_clk,                                          --            clock.clk
			wb_rst_i   => rst_controller_001_reset_out_reset,                         --            reset.reset
			wb_inta_o  => irq_mapper_002_receiver2_irq                                -- interrupt_sender.irq
		);

	i2c_master_is2 : component i2c_opencores
		port map (
			wb_adr_i   => mm_interconnect_0_i2c_master_is2_avalon_slave_0_address,    --   avalon_slave_0.address
			wb_dat_i   => mm_interconnect_0_i2c_master_is2_avalon_slave_0_writedata,  --                 .writedata
			wb_dat_o   => mm_interconnect_0_i2c_master_is2_avalon_slave_0_readdata,   --                 .readdata
			wb_we_i    => mm_interconnect_0_i2c_master_is2_avalon_slave_0_write,      --                 .write
			wb_stb_i   => mm_interconnect_0_i2c_master_is2_avalon_slave_0_chipselect, --                 .chipselect
			wb_ack_o   => i2c_master_is2_avalon_slave_0_waitrequest,                  --                 .waitrequest_n
			scl_pad_io => i2c_master_is2_conduit_end_scl,                             --      conduit_end.scl
			sda_pad_io => i2c_master_is2_conduit_end_sda,                             --                 .sda
			wb_clk_i   => pll_0_outclk0_clk,                                          --            clock.clk
			wb_rst_i   => rst_controller_001_reset_out_reset,                         --            reset.reset
			wb_inta_o  => irq_mapper_002_receiver3_irq                                -- interrupt_sender.irq
		);

	i2c_master_is3 : component i2c_opencores
		port map (
			wb_adr_i   => mm_interconnect_0_i2c_master_is3_avalon_slave_0_address,    --   avalon_slave_0.address
			wb_dat_i   => mm_interconnect_0_i2c_master_is3_avalon_slave_0_writedata,  --                 .writedata
			wb_dat_o   => mm_interconnect_0_i2c_master_is3_avalon_slave_0_readdata,   --                 .readdata
			wb_we_i    => mm_interconnect_0_i2c_master_is3_avalon_slave_0_write,      --                 .write
			wb_stb_i   => mm_interconnect_0_i2c_master_is3_avalon_slave_0_chipselect, --                 .chipselect
			wb_ack_o   => i2c_master_is3_avalon_slave_0_waitrequest,                  --                 .waitrequest_n
			scl_pad_io => i2c_master_is3_conduit_end_scl,                             --      conduit_end.scl
			sda_pad_io => i2c_master_is3_conduit_end_sda,                             --                 .sda
			wb_clk_i   => pll_0_outclk0_clk,                                          --            clock.clk
			wb_rst_i   => rst_controller_001_reset_out_reset,                         --            reset.reset
			wb_inta_o  => irq_mapper_002_receiver4_irq                                -- interrupt_sender.irq
		);

	i2c_master_is4 : component i2c_opencores
		port map (
			wb_adr_i   => mm_interconnect_0_i2c_master_is4_avalon_slave_0_address,    --   avalon_slave_0.address
			wb_dat_i   => mm_interconnect_0_i2c_master_is4_avalon_slave_0_writedata,  --                 .writedata
			wb_dat_o   => mm_interconnect_0_i2c_master_is4_avalon_slave_0_readdata,   --                 .readdata
			wb_we_i    => mm_interconnect_0_i2c_master_is4_avalon_slave_0_write,      --                 .write
			wb_stb_i   => mm_interconnect_0_i2c_master_is4_avalon_slave_0_chipselect, --                 .chipselect
			wb_ack_o   => i2c_master_is4_avalon_slave_0_waitrequest,                  --                 .waitrequest_n
			scl_pad_io => i2c_master_is4_conduit_end_scl,                             --      conduit_end.scl
			sda_pad_io => i2c_master_is4_conduit_end_sda,                             --                 .sda
			wb_clk_i   => pll_0_outclk0_clk,                                          --            clock.clk
			wb_rst_i   => rst_controller_001_reset_out_reset,                         --            reset.reset
			wb_inta_o  => irq_mapper_002_receiver5_irq                                -- interrupt_sender.irq
		);

	onchip_memory_nios_cpu : component fluid_board_soc_onchip_memory_nios_cpu
		port map (
			address     => mm_interconnect_0_onchip_memory_nios_cpu_s1_address,    --     s1.address
			clken       => mm_interconnect_0_onchip_memory_nios_cpu_s1_clken,      --       .clken
			chipselect  => mm_interconnect_0_onchip_memory_nios_cpu_s1_chipselect, --       .chipselect
			write       => mm_interconnect_0_onchip_memory_nios_cpu_s1_write,      --       .write
			readdata    => mm_interconnect_0_onchip_memory_nios_cpu_s1_readdata,   --       .readdata
			writedata   => mm_interconnect_0_onchip_memory_nios_cpu_s1_writedata,  --       .writedata
			byteenable  => mm_interconnect_0_onchip_memory_nios_cpu_s1_byteenable, --       .byteenable
			address2    => mm_interconnect_1_onchip_memory_nios_cpu_s2_address,    --     s2.address
			chipselect2 => mm_interconnect_1_onchip_memory_nios_cpu_s2_chipselect, --       .chipselect
			clken2      => mm_interconnect_1_onchip_memory_nios_cpu_s2_clken,      --       .clken
			write2      => mm_interconnect_1_onchip_memory_nios_cpu_s2_write,      --       .write
			readdata2   => mm_interconnect_1_onchip_memory_nios_cpu_s2_readdata,   --       .readdata
			writedata2  => mm_interconnect_1_onchip_memory_nios_cpu_s2_writedata,  --       .writedata
			byteenable2 => mm_interconnect_1_onchip_memory_nios_cpu_s2_byteenable, --       .byteenable
			clk         => pll_0_outclk0_clk,                                      --   clk1.clk
			reset       => rst_controller_reset_out_reset,                         -- reset1.reset
			reset_req   => rst_controller_reset_out_reset_req                      --       .reset_req
		);

	pio_input : component fluid_board_soc_pio_input
		port map (
			clk        => pll_0_outclk0_clk,                              --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_pio_input_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_input_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_input_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_input_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_input_s1_readdata,        --                    .readdata
			in_port    => pio_input_external_connection_export,           -- external_connection.export
			irq        => irq_mapper_002_receiver6_irq                    --                 irq.irq
		);

	pio_output : component fluid_board_soc_pio_output
		port map (
			clk        => pll_0_outclk0_clk,                               --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_0_pio_output_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_output_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_output_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_output_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_output_s1_readdata,        --                    .readdata
			out_port   => pio_output_external_connection_export            -- external_connection.export
		);

	onchip_memory_nios_arm : component fluid_board_soc_onchip_memory_nios_arm
		port map (
			address     => mm_interconnect_0_onchip_memory_nios_arm_s1_address,    --     s1.address
			clken       => mm_interconnect_0_onchip_memory_nios_arm_s1_clken,      --       .clken
			chipselect  => mm_interconnect_0_onchip_memory_nios_arm_s1_chipselect, --       .chipselect
			write       => mm_interconnect_0_onchip_memory_nios_arm_s1_write,      --       .write
			readdata    => mm_interconnect_0_onchip_memory_nios_arm_s1_readdata,   --       .readdata
			writedata   => mm_interconnect_0_onchip_memory_nios_arm_s1_writedata,  --       .writedata
			byteenable  => mm_interconnect_0_onchip_memory_nios_arm_s1_byteenable, --       .byteenable
			address2    => mm_interconnect_1_onchip_memory_nios_arm_s2_address,    --     s2.address
			chipselect2 => mm_interconnect_1_onchip_memory_nios_arm_s2_chipselect, --       .chipselect
			clken2      => mm_interconnect_1_onchip_memory_nios_arm_s2_clken,      --       .clken
			write2      => mm_interconnect_1_onchip_memory_nios_arm_s2_write,      --       .write
			readdata2   => mm_interconnect_1_onchip_memory_nios_arm_s2_readdata,   --       .readdata
			writedata2  => mm_interconnect_1_onchip_memory_nios_arm_s2_writedata,  --       .writedata
			byteenable2 => mm_interconnect_1_onchip_memory_nios_arm_s2_byteenable, --       .byteenable
			clk         => pll_0_outclk0_clk,                                      --   clk1.clk
			reset       => rst_controller_reset_out_reset,                         -- reset1.reset
			reset_req   => rst_controller_reset_out_reset_req                      --       .reset_req
		);

	jtag_uart : component fluid_board_soc_jtag_uart
		port map (
			clk            => pll_0_outclk0_clk,                                             --               clk.clk
			rst_n          => rst_controller_001_reset_out_reset_ports_inv,                  --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                       --               irq.irq
		);

	fpga_only_master : component fluid_board_soc_fpga_only_master
		port map (
			clk_clk              => pll_0_outclk0_clk,                     --          clk.clk
			clk_reset_reset      => qsys_reset_reset_n_ports_inv,          --    clk_reset.reset
			master_address       => fpga_only_master_master_address,       --       master.address
			master_readdata      => fpga_only_master_master_readdata,      --             .readdata
			master_read          => fpga_only_master_master_read,          --             .read
			master_write         => fpga_only_master_master_write,         --             .write
			master_writedata     => fpga_only_master_master_writedata,     --             .writedata
			master_waitrequest   => fpga_only_master_master_waitrequest,   --             .waitrequest
			master_readdatavalid => fpga_only_master_master_readdatavalid, --             .readdatavalid
			master_byteenable    => fpga_only_master_master_byteenable,    --             .byteenable
			master_reset_reset   => open                                   -- master_reset.reset
		);

	i2c_master_d : component i2c_opencores
		port map (
			wb_adr_i   => mm_interconnect_0_i2c_master_d_avalon_slave_0_address,    --   avalon_slave_0.address
			wb_dat_i   => mm_interconnect_0_i2c_master_d_avalon_slave_0_writedata,  --                 .writedata
			wb_dat_o   => mm_interconnect_0_i2c_master_d_avalon_slave_0_readdata,   --                 .readdata
			wb_we_i    => mm_interconnect_0_i2c_master_d_avalon_slave_0_write,      --                 .write
			wb_stb_i   => mm_interconnect_0_i2c_master_d_avalon_slave_0_chipselect, --                 .chipselect
			wb_ack_o   => i2c_master_d_avalon_slave_0_waitrequest,                  --                 .waitrequest_n
			scl_pad_io => i2c_master_d_conduit_end_scl,                             --      conduit_end.scl
			sda_pad_io => i2c_master_d_conduit_end_sda,                             --                 .sda
			wb_clk_i   => pll_0_outclk0_clk,                                        --            clock.clk
			wb_rst_i   => rst_controller_001_reset_out_reset,                       --            reset.reset
			wb_inta_o  => irq_mapper_002_receiver8_irq                              -- interrupt_sender.irq
		);

	i2c_master_f : component i2c_opencores
		port map (
			wb_adr_i   => mm_interconnect_0_i2c_master_f_avalon_slave_0_address,    --   avalon_slave_0.address
			wb_dat_i   => mm_interconnect_0_i2c_master_f_avalon_slave_0_writedata,  --                 .writedata
			wb_dat_o   => mm_interconnect_0_i2c_master_f_avalon_slave_0_readdata,   --                 .readdata
			wb_we_i    => mm_interconnect_0_i2c_master_f_avalon_slave_0_write,      --                 .write
			wb_stb_i   => mm_interconnect_0_i2c_master_f_avalon_slave_0_chipselect, --                 .chipselect
			wb_ack_o   => i2c_master_f_avalon_slave_0_waitrequest,                  --                 .waitrequest_n
			scl_pad_io => i2c_master_f_conduit_end_scl,                             --      conduit_end.scl
			sda_pad_io => i2c_master_f_conduit_end_sda,                             --                 .sda
			wb_clk_i   => pll_0_outclk0_clk,                                        --            clock.clk
			wb_rst_i   => rst_controller_001_reset_out_reset,                       --            reset.reset
			wb_inta_o  => irq_mapper_002_receiver9_irq                              -- interrupt_sender.irq
		);

	i2c_master_p : component i2c_opencores
		port map (
			wb_adr_i   => mm_interconnect_0_i2c_master_p_avalon_slave_0_address,    --   avalon_slave_0.address
			wb_dat_i   => mm_interconnect_0_i2c_master_p_avalon_slave_0_writedata,  --                 .writedata
			wb_dat_o   => mm_interconnect_0_i2c_master_p_avalon_slave_0_readdata,   --                 .readdata
			wb_we_i    => mm_interconnect_0_i2c_master_p_avalon_slave_0_write,      --                 .write
			wb_stb_i   => mm_interconnect_0_i2c_master_p_avalon_slave_0_chipselect, --                 .chipselect
			wb_ack_o   => i2c_master_p_avalon_slave_0_waitrequest,                  --                 .waitrequest_n
			scl_pad_io => i2c_master_p_conduit_end_scl,                             --      conduit_end.scl
			sda_pad_io => i2c_master_p_conduit_end_sda,                             --                 .sda
			wb_clk_i   => pll_0_outclk0_clk,                                        --            clock.clk
			wb_rst_i   => rst_controller_001_reset_out_reset,                       --            reset.reset
			wb_inta_o  => irq_mapper_002_receiver10_irq                             -- interrupt_sender.irq
		);

	pio_reset_nios : component fluid_board_soc_pio_reset_nios
		port map (
			clk        => pll_0_outclk0_clk,                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,            --               reset.reset_n
			address    => mm_interconnect_0_pio_reset_nios_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_reset_nios_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_reset_nios_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_reset_nios_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_reset_nios_s1_readdata,        --                    .readdata
			out_port   => pio_reset_nios_external_connection_export            -- external_connection.export
		);

	mm_interconnect_0 : component fluid_board_soc_mm_interconnect_0
		port map (
			hps_0_h2f_lw_axi_master_awid                                        => hps_0_h2f_lw_axi_master_awid,                                 --                                       hps_0_h2f_lw_axi_master.awid
			hps_0_h2f_lw_axi_master_awaddr                                      => hps_0_h2f_lw_axi_master_awaddr,                               --                                                              .awaddr
			hps_0_h2f_lw_axi_master_awlen                                       => hps_0_h2f_lw_axi_master_awlen,                                --                                                              .awlen
			hps_0_h2f_lw_axi_master_awsize                                      => hps_0_h2f_lw_axi_master_awsize,                               --                                                              .awsize
			hps_0_h2f_lw_axi_master_awburst                                     => hps_0_h2f_lw_axi_master_awburst,                              --                                                              .awburst
			hps_0_h2f_lw_axi_master_awlock                                      => hps_0_h2f_lw_axi_master_awlock,                               --                                                              .awlock
			hps_0_h2f_lw_axi_master_awcache                                     => hps_0_h2f_lw_axi_master_awcache,                              --                                                              .awcache
			hps_0_h2f_lw_axi_master_awprot                                      => hps_0_h2f_lw_axi_master_awprot,                               --                                                              .awprot
			hps_0_h2f_lw_axi_master_awvalid                                     => hps_0_h2f_lw_axi_master_awvalid,                              --                                                              .awvalid
			hps_0_h2f_lw_axi_master_awready                                     => hps_0_h2f_lw_axi_master_awready,                              --                                                              .awready
			hps_0_h2f_lw_axi_master_wid                                         => hps_0_h2f_lw_axi_master_wid,                                  --                                                              .wid
			hps_0_h2f_lw_axi_master_wdata                                       => hps_0_h2f_lw_axi_master_wdata,                                --                                                              .wdata
			hps_0_h2f_lw_axi_master_wstrb                                       => hps_0_h2f_lw_axi_master_wstrb,                                --                                                              .wstrb
			hps_0_h2f_lw_axi_master_wlast                                       => hps_0_h2f_lw_axi_master_wlast,                                --                                                              .wlast
			hps_0_h2f_lw_axi_master_wvalid                                      => hps_0_h2f_lw_axi_master_wvalid,                               --                                                              .wvalid
			hps_0_h2f_lw_axi_master_wready                                      => hps_0_h2f_lw_axi_master_wready,                               --                                                              .wready
			hps_0_h2f_lw_axi_master_bid                                         => hps_0_h2f_lw_axi_master_bid,                                  --                                                              .bid
			hps_0_h2f_lw_axi_master_bresp                                       => hps_0_h2f_lw_axi_master_bresp,                                --                                                              .bresp
			hps_0_h2f_lw_axi_master_bvalid                                      => hps_0_h2f_lw_axi_master_bvalid,                               --                                                              .bvalid
			hps_0_h2f_lw_axi_master_bready                                      => hps_0_h2f_lw_axi_master_bready,                               --                                                              .bready
			hps_0_h2f_lw_axi_master_arid                                        => hps_0_h2f_lw_axi_master_arid,                                 --                                                              .arid
			hps_0_h2f_lw_axi_master_araddr                                      => hps_0_h2f_lw_axi_master_araddr,                               --                                                              .araddr
			hps_0_h2f_lw_axi_master_arlen                                       => hps_0_h2f_lw_axi_master_arlen,                                --                                                              .arlen
			hps_0_h2f_lw_axi_master_arsize                                      => hps_0_h2f_lw_axi_master_arsize,                               --                                                              .arsize
			hps_0_h2f_lw_axi_master_arburst                                     => hps_0_h2f_lw_axi_master_arburst,                              --                                                              .arburst
			hps_0_h2f_lw_axi_master_arlock                                      => hps_0_h2f_lw_axi_master_arlock,                               --                                                              .arlock
			hps_0_h2f_lw_axi_master_arcache                                     => hps_0_h2f_lw_axi_master_arcache,                              --                                                              .arcache
			hps_0_h2f_lw_axi_master_arprot                                      => hps_0_h2f_lw_axi_master_arprot,                               --                                                              .arprot
			hps_0_h2f_lw_axi_master_arvalid                                     => hps_0_h2f_lw_axi_master_arvalid,                              --                                                              .arvalid
			hps_0_h2f_lw_axi_master_arready                                     => hps_0_h2f_lw_axi_master_arready,                              --                                                              .arready
			hps_0_h2f_lw_axi_master_rid                                         => hps_0_h2f_lw_axi_master_rid,                                  --                                                              .rid
			hps_0_h2f_lw_axi_master_rdata                                       => hps_0_h2f_lw_axi_master_rdata,                                --                                                              .rdata
			hps_0_h2f_lw_axi_master_rresp                                       => hps_0_h2f_lw_axi_master_rresp,                                --                                                              .rresp
			hps_0_h2f_lw_axi_master_rlast                                       => hps_0_h2f_lw_axi_master_rlast,                                --                                                              .rlast
			hps_0_h2f_lw_axi_master_rvalid                                      => hps_0_h2f_lw_axi_master_rvalid,                               --                                                              .rvalid
			hps_0_h2f_lw_axi_master_rready                                      => hps_0_h2f_lw_axi_master_rready,                               --                                                              .rready
			clk_i_clk_clk                                                       => pll_0_outclk0_clk,                                            --                                                     clk_i_clk.clk
			fpga_only_master_clk_reset_reset_bridge_in_reset_reset              => rst_controller_001_reset_out_reset,                           --              fpga_only_master_clk_reset_reset_bridge_in_reset.reset
			hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset => rst_controller_002_reset_out_reset,                           -- hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
			nios2_qsys_0_reset_n_reset_bridge_in_reset_reset                    => rst_controller_001_reset_out_reset,                           --                    nios2_qsys_0_reset_n_reset_bridge_in_reset.reset
			sysid_reset_reset_bridge_in_reset_reset                             => rst_controller_reset_out_reset,                               --                             sysid_reset_reset_bridge_in_reset.reset
			fpga_only_master_master_address                                     => fpga_only_master_master_address,                              --                                       fpga_only_master_master.address
			fpga_only_master_master_waitrequest                                 => fpga_only_master_master_waitrequest,                          --                                                              .waitrequest
			fpga_only_master_master_byteenable                                  => fpga_only_master_master_byteenable,                           --                                                              .byteenable
			fpga_only_master_master_read                                        => fpga_only_master_master_read,                                 --                                                              .read
			fpga_only_master_master_readdata                                    => fpga_only_master_master_readdata,                             --                                                              .readdata
			fpga_only_master_master_readdatavalid                               => fpga_only_master_master_readdatavalid,                        --                                                              .readdatavalid
			fpga_only_master_master_write                                       => fpga_only_master_master_write,                                --                                                              .write
			fpga_only_master_master_writedata                                   => fpga_only_master_master_writedata,                            --                                                              .writedata
			nios2_qsys_0_data_master_address                                    => nios2_qsys_0_data_master_address,                             --                                      nios2_qsys_0_data_master.address
			nios2_qsys_0_data_master_waitrequest                                => nios2_qsys_0_data_master_waitrequest,                         --                                                              .waitrequest
			nios2_qsys_0_data_master_byteenable                                 => nios2_qsys_0_data_master_byteenable,                          --                                                              .byteenable
			nios2_qsys_0_data_master_read                                       => nios2_qsys_0_data_master_read,                                --                                                              .read
			nios2_qsys_0_data_master_readdata                                   => nios2_qsys_0_data_master_readdata,                            --                                                              .readdata
			nios2_qsys_0_data_master_write                                      => nios2_qsys_0_data_master_write,                               --                                                              .write
			nios2_qsys_0_data_master_writedata                                  => nios2_qsys_0_data_master_writedata,                           --                                                              .writedata
			nios2_qsys_0_data_master_debugaccess                                => nios2_qsys_0_data_master_debugaccess,                         --                                                              .debugaccess
			nios2_qsys_0_instruction_master_address                             => nios2_qsys_0_instruction_master_address,                      --                               nios2_qsys_0_instruction_master.address
			nios2_qsys_0_instruction_master_waitrequest                         => nios2_qsys_0_instruction_master_waitrequest,                  --                                                              .waitrequest
			nios2_qsys_0_instruction_master_read                                => nios2_qsys_0_instruction_master_read,                         --                                                              .read
			nios2_qsys_0_instruction_master_readdata                            => nios2_qsys_0_instruction_master_readdata,                     --                                                              .readdata
			nios2_qsys_0_instruction_master_readdatavalid                       => nios2_qsys_0_instruction_master_readdatavalid,                --                                                              .readdatavalid
			avalon_spi_AMC7891_0_s1_address                                     => mm_interconnect_0_avalon_spi_amc7891_0_s1_address,            --                                       avalon_spi_AMC7891_0_s1.address
			avalon_spi_AMC7891_0_s1_write                                       => mm_interconnect_0_avalon_spi_amc7891_0_s1_write,              --                                                              .write
			avalon_spi_AMC7891_0_s1_read                                        => mm_interconnect_0_avalon_spi_amc7891_0_s1_read,               --                                                              .read
			avalon_spi_AMC7891_0_s1_readdata                                    => mm_interconnect_0_avalon_spi_amc7891_0_s1_readdata,           --                                                              .readdata
			avalon_spi_AMC7891_0_s1_writedata                                   => mm_interconnect_0_avalon_spi_amc7891_0_s1_writedata,          --                                                              .writedata
			avalon_spi_AMC7891_0_s1_waitrequest                                 => mm_interconnect_0_avalon_spi_amc7891_0_s1_waitrequest,        --                                                              .waitrequest
			avalon_spi_AMC7891_1_s1_address                                     => mm_interconnect_0_avalon_spi_amc7891_1_s1_address,            --                                       avalon_spi_AMC7891_1_s1.address
			avalon_spi_AMC7891_1_s1_write                                       => mm_interconnect_0_avalon_spi_amc7891_1_s1_write,              --                                                              .write
			avalon_spi_AMC7891_1_s1_read                                        => mm_interconnect_0_avalon_spi_amc7891_1_s1_read,               --                                                              .read
			avalon_spi_AMC7891_1_s1_readdata                                    => mm_interconnect_0_avalon_spi_amc7891_1_s1_readdata,           --                                                              .readdata
			avalon_spi_AMC7891_1_s1_writedata                                   => mm_interconnect_0_avalon_spi_amc7891_1_s1_writedata,          --                                                              .writedata
			avalon_spi_AMC7891_1_s1_waitrequest                                 => mm_interconnect_0_avalon_spi_amc7891_1_s1_waitrequest,        --                                                              .waitrequest
			i2c_master_d_avalon_slave_0_address                                 => mm_interconnect_0_i2c_master_d_avalon_slave_0_address,        --                                   i2c_master_d_avalon_slave_0.address
			i2c_master_d_avalon_slave_0_write                                   => mm_interconnect_0_i2c_master_d_avalon_slave_0_write,          --                                                              .write
			i2c_master_d_avalon_slave_0_readdata                                => mm_interconnect_0_i2c_master_d_avalon_slave_0_readdata,       --                                                              .readdata
			i2c_master_d_avalon_slave_0_writedata                               => mm_interconnect_0_i2c_master_d_avalon_slave_0_writedata,      --                                                              .writedata
			i2c_master_d_avalon_slave_0_waitrequest                             => mm_interconnect_0_i2c_master_d_avalon_slave_0_inv,            --                                                              .waitrequest
			i2c_master_d_avalon_slave_0_chipselect                              => mm_interconnect_0_i2c_master_d_avalon_slave_0_chipselect,     --                                                              .chipselect
			i2c_master_f_avalon_slave_0_address                                 => mm_interconnect_0_i2c_master_f_avalon_slave_0_address,        --                                   i2c_master_f_avalon_slave_0.address
			i2c_master_f_avalon_slave_0_write                                   => mm_interconnect_0_i2c_master_f_avalon_slave_0_write,          --                                                              .write
			i2c_master_f_avalon_slave_0_readdata                                => mm_interconnect_0_i2c_master_f_avalon_slave_0_readdata,       --                                                              .readdata
			i2c_master_f_avalon_slave_0_writedata                               => mm_interconnect_0_i2c_master_f_avalon_slave_0_writedata,      --                                                              .writedata
			i2c_master_f_avalon_slave_0_waitrequest                             => mm_interconnect_0_i2c_master_f_avalon_slave_0_inv,            --                                                              .waitrequest
			i2c_master_f_avalon_slave_0_chipselect                              => mm_interconnect_0_i2c_master_f_avalon_slave_0_chipselect,     --                                                              .chipselect
			i2c_master_is1_avalon_slave_0_address                               => mm_interconnect_0_i2c_master_is1_avalon_slave_0_address,      --                                 i2c_master_is1_avalon_slave_0.address
			i2c_master_is1_avalon_slave_0_write                                 => mm_interconnect_0_i2c_master_is1_avalon_slave_0_write,        --                                                              .write
			i2c_master_is1_avalon_slave_0_readdata                              => mm_interconnect_0_i2c_master_is1_avalon_slave_0_readdata,     --                                                              .readdata
			i2c_master_is1_avalon_slave_0_writedata                             => mm_interconnect_0_i2c_master_is1_avalon_slave_0_writedata,    --                                                              .writedata
			i2c_master_is1_avalon_slave_0_waitrequest                           => mm_interconnect_0_i2c_master_is1_avalon_slave_0_inv,          --                                                              .waitrequest
			i2c_master_is1_avalon_slave_0_chipselect                            => mm_interconnect_0_i2c_master_is1_avalon_slave_0_chipselect,   --                                                              .chipselect
			i2c_master_is2_avalon_slave_0_address                               => mm_interconnect_0_i2c_master_is2_avalon_slave_0_address,      --                                 i2c_master_is2_avalon_slave_0.address
			i2c_master_is2_avalon_slave_0_write                                 => mm_interconnect_0_i2c_master_is2_avalon_slave_0_write,        --                                                              .write
			i2c_master_is2_avalon_slave_0_readdata                              => mm_interconnect_0_i2c_master_is2_avalon_slave_0_readdata,     --                                                              .readdata
			i2c_master_is2_avalon_slave_0_writedata                             => mm_interconnect_0_i2c_master_is2_avalon_slave_0_writedata,    --                                                              .writedata
			i2c_master_is2_avalon_slave_0_waitrequest                           => mm_interconnect_0_i2c_master_is2_avalon_slave_0_inv,          --                                                              .waitrequest
			i2c_master_is2_avalon_slave_0_chipselect                            => mm_interconnect_0_i2c_master_is2_avalon_slave_0_chipselect,   --                                                              .chipselect
			i2c_master_is3_avalon_slave_0_address                               => mm_interconnect_0_i2c_master_is3_avalon_slave_0_address,      --                                 i2c_master_is3_avalon_slave_0.address
			i2c_master_is3_avalon_slave_0_write                                 => mm_interconnect_0_i2c_master_is3_avalon_slave_0_write,        --                                                              .write
			i2c_master_is3_avalon_slave_0_readdata                              => mm_interconnect_0_i2c_master_is3_avalon_slave_0_readdata,     --                                                              .readdata
			i2c_master_is3_avalon_slave_0_writedata                             => mm_interconnect_0_i2c_master_is3_avalon_slave_0_writedata,    --                                                              .writedata
			i2c_master_is3_avalon_slave_0_waitrequest                           => mm_interconnect_0_i2c_master_is3_avalon_slave_0_inv,          --                                                              .waitrequest
			i2c_master_is3_avalon_slave_0_chipselect                            => mm_interconnect_0_i2c_master_is3_avalon_slave_0_chipselect,   --                                                              .chipselect
			i2c_master_is4_avalon_slave_0_address                               => mm_interconnect_0_i2c_master_is4_avalon_slave_0_address,      --                                 i2c_master_is4_avalon_slave_0.address
			i2c_master_is4_avalon_slave_0_write                                 => mm_interconnect_0_i2c_master_is4_avalon_slave_0_write,        --                                                              .write
			i2c_master_is4_avalon_slave_0_readdata                              => mm_interconnect_0_i2c_master_is4_avalon_slave_0_readdata,     --                                                              .readdata
			i2c_master_is4_avalon_slave_0_writedata                             => mm_interconnect_0_i2c_master_is4_avalon_slave_0_writedata,    --                                                              .writedata
			i2c_master_is4_avalon_slave_0_waitrequest                           => mm_interconnect_0_i2c_master_is4_avalon_slave_0_inv,          --                                                              .waitrequest
			i2c_master_is4_avalon_slave_0_chipselect                            => mm_interconnect_0_i2c_master_is4_avalon_slave_0_chipselect,   --                                                              .chipselect
			i2c_master_p_avalon_slave_0_address                                 => mm_interconnect_0_i2c_master_p_avalon_slave_0_address,        --                                   i2c_master_p_avalon_slave_0.address
			i2c_master_p_avalon_slave_0_write                                   => mm_interconnect_0_i2c_master_p_avalon_slave_0_write,          --                                                              .write
			i2c_master_p_avalon_slave_0_readdata                                => mm_interconnect_0_i2c_master_p_avalon_slave_0_readdata,       --                                                              .readdata
			i2c_master_p_avalon_slave_0_writedata                               => mm_interconnect_0_i2c_master_p_avalon_slave_0_writedata,      --                                                              .writedata
			i2c_master_p_avalon_slave_0_waitrequest                             => mm_interconnect_0_i2c_master_p_avalon_slave_0_inv,            --                                                              .waitrequest
			i2c_master_p_avalon_slave_0_chipselect                              => mm_interconnect_0_i2c_master_p_avalon_slave_0_chipselect,     --                                                              .chipselect
			jtag_uart_avalon_jtag_slave_address                                 => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,        --                                   jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write                                   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,          --                                                              .write
			jtag_uart_avalon_jtag_slave_read                                    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,           --                                                              .read
			jtag_uart_avalon_jtag_slave_readdata                                => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,       --                                                              .readdata
			jtag_uart_avalon_jtag_slave_writedata                               => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,      --                                                              .writedata
			jtag_uart_avalon_jtag_slave_waitrequest                             => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,    --                                                              .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                              => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,     --                                                              .chipselect
			nios2_qsys_0_jtag_debug_module_address                              => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address,     --                                nios2_qsys_0_jtag_debug_module.address
			nios2_qsys_0_jtag_debug_module_write                                => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write,       --                                                              .write
			nios2_qsys_0_jtag_debug_module_read                                 => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read,        --                                                              .read
			nios2_qsys_0_jtag_debug_module_readdata                             => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata,    --                                                              .readdata
			nios2_qsys_0_jtag_debug_module_writedata                            => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata,   --                                                              .writedata
			nios2_qsys_0_jtag_debug_module_byteenable                           => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable,  --                                                              .byteenable
			nios2_qsys_0_jtag_debug_module_waitrequest                          => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest, --                                                              .waitrequest
			nios2_qsys_0_jtag_debug_module_debugaccess                          => mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess, --                                                              .debugaccess
			onchip_memory_nios_arm_s1_address                                   => mm_interconnect_0_onchip_memory_nios_arm_s1_address,          --                                     onchip_memory_nios_arm_s1.address
			onchip_memory_nios_arm_s1_write                                     => mm_interconnect_0_onchip_memory_nios_arm_s1_write,            --                                                              .write
			onchip_memory_nios_arm_s1_readdata                                  => mm_interconnect_0_onchip_memory_nios_arm_s1_readdata,         --                                                              .readdata
			onchip_memory_nios_arm_s1_writedata                                 => mm_interconnect_0_onchip_memory_nios_arm_s1_writedata,        --                                                              .writedata
			onchip_memory_nios_arm_s1_byteenable                                => mm_interconnect_0_onchip_memory_nios_arm_s1_byteenable,       --                                                              .byteenable
			onchip_memory_nios_arm_s1_chipselect                                => mm_interconnect_0_onchip_memory_nios_arm_s1_chipselect,       --                                                              .chipselect
			onchip_memory_nios_arm_s1_clken                                     => mm_interconnect_0_onchip_memory_nios_arm_s1_clken,            --                                                              .clken
			onchip_memory_nios_cpu_s1_address                                   => mm_interconnect_0_onchip_memory_nios_cpu_s1_address,          --                                     onchip_memory_nios_cpu_s1.address
			onchip_memory_nios_cpu_s1_write                                     => mm_interconnect_0_onchip_memory_nios_cpu_s1_write,            --                                                              .write
			onchip_memory_nios_cpu_s1_readdata                                  => mm_interconnect_0_onchip_memory_nios_cpu_s1_readdata,         --                                                              .readdata
			onchip_memory_nios_cpu_s1_writedata                                 => mm_interconnect_0_onchip_memory_nios_cpu_s1_writedata,        --                                                              .writedata
			onchip_memory_nios_cpu_s1_byteenable                                => mm_interconnect_0_onchip_memory_nios_cpu_s1_byteenable,       --                                                              .byteenable
			onchip_memory_nios_cpu_s1_chipselect                                => mm_interconnect_0_onchip_memory_nios_cpu_s1_chipselect,       --                                                              .chipselect
			onchip_memory_nios_cpu_s1_clken                                     => mm_interconnect_0_onchip_memory_nios_cpu_s1_clken,            --                                                              .clken
			pio_input_s1_address                                                => mm_interconnect_0_pio_input_s1_address,                       --                                                  pio_input_s1.address
			pio_input_s1_write                                                  => mm_interconnect_0_pio_input_s1_write,                         --                                                              .write
			pio_input_s1_readdata                                               => mm_interconnect_0_pio_input_s1_readdata,                      --                                                              .readdata
			pio_input_s1_writedata                                              => mm_interconnect_0_pio_input_s1_writedata,                     --                                                              .writedata
			pio_input_s1_chipselect                                             => mm_interconnect_0_pio_input_s1_chipselect,                    --                                                              .chipselect
			pio_output_s1_address                                               => mm_interconnect_0_pio_output_s1_address,                      --                                                 pio_output_s1.address
			pio_output_s1_write                                                 => mm_interconnect_0_pio_output_s1_write,                        --                                                              .write
			pio_output_s1_readdata                                              => mm_interconnect_0_pio_output_s1_readdata,                     --                                                              .readdata
			pio_output_s1_writedata                                             => mm_interconnect_0_pio_output_s1_writedata,                    --                                                              .writedata
			pio_output_s1_chipselect                                            => mm_interconnect_0_pio_output_s1_chipselect,                   --                                                              .chipselect
			pio_reset_nios_s1_address                                           => mm_interconnect_0_pio_reset_nios_s1_address,                  --                                             pio_reset_nios_s1.address
			pio_reset_nios_s1_write                                             => mm_interconnect_0_pio_reset_nios_s1_write,                    --                                                              .write
			pio_reset_nios_s1_readdata                                          => mm_interconnect_0_pio_reset_nios_s1_readdata,                 --                                                              .readdata
			pio_reset_nios_s1_writedata                                         => mm_interconnect_0_pio_reset_nios_s1_writedata,                --                                                              .writedata
			pio_reset_nios_s1_chipselect                                        => mm_interconnect_0_pio_reset_nios_s1_chipselect,               --                                                              .chipselect
			sysid_control_slave_address                                         => mm_interconnect_0_sysid_control_slave_address,                --                                           sysid_control_slave.address
			sysid_control_slave_readdata                                        => mm_interconnect_0_sysid_control_slave_readdata,               --                                                              .readdata
			timer_0_s1_address                                                  => mm_interconnect_0_timer_0_s1_address,                         --                                                    timer_0_s1.address
			timer_0_s1_write                                                    => mm_interconnect_0_timer_0_s1_write,                           --                                                              .write
			timer_0_s1_readdata                                                 => mm_interconnect_0_timer_0_s1_readdata,                        --                                                              .readdata
			timer_0_s1_writedata                                                => mm_interconnect_0_timer_0_s1_writedata,                       --                                                              .writedata
			timer_0_s1_chipselect                                               => mm_interconnect_0_timer_0_s1_chipselect,                      --                                                              .chipselect
			timer_1_s1_address                                                  => mm_interconnect_0_timer_1_s1_address,                         --                                                    timer_1_s1.address
			timer_1_s1_write                                                    => mm_interconnect_0_timer_1_s1_write,                           --                                                              .write
			timer_1_s1_readdata                                                 => mm_interconnect_0_timer_1_s1_readdata,                        --                                                              .readdata
			timer_1_s1_writedata                                                => mm_interconnect_0_timer_1_s1_writedata,                       --                                                              .writedata
			timer_1_s1_chipselect                                               => mm_interconnect_0_timer_1_s1_chipselect                       --                                                              .chipselect
		);

	mm_interconnect_1 : component fluid_board_soc_mm_interconnect_1
		port map (
			hps_0_h2f_axi_master_awid                                        => hps_0_h2f_axi_master_awid,                                      --                                       hps_0_h2f_axi_master.awid
			hps_0_h2f_axi_master_awaddr                                      => hps_0_h2f_axi_master_awaddr,                                    --                                                           .awaddr
			hps_0_h2f_axi_master_awlen                                       => hps_0_h2f_axi_master_awlen,                                     --                                                           .awlen
			hps_0_h2f_axi_master_awsize                                      => hps_0_h2f_axi_master_awsize,                                    --                                                           .awsize
			hps_0_h2f_axi_master_awburst                                     => hps_0_h2f_axi_master_awburst,                                   --                                                           .awburst
			hps_0_h2f_axi_master_awlock                                      => hps_0_h2f_axi_master_awlock,                                    --                                                           .awlock
			hps_0_h2f_axi_master_awcache                                     => hps_0_h2f_axi_master_awcache,                                   --                                                           .awcache
			hps_0_h2f_axi_master_awprot                                      => hps_0_h2f_axi_master_awprot,                                    --                                                           .awprot
			hps_0_h2f_axi_master_awvalid                                     => hps_0_h2f_axi_master_awvalid,                                   --                                                           .awvalid
			hps_0_h2f_axi_master_awready                                     => hps_0_h2f_axi_master_awready,                                   --                                                           .awready
			hps_0_h2f_axi_master_wid                                         => hps_0_h2f_axi_master_wid,                                       --                                                           .wid
			hps_0_h2f_axi_master_wdata                                       => hps_0_h2f_axi_master_wdata,                                     --                                                           .wdata
			hps_0_h2f_axi_master_wstrb                                       => hps_0_h2f_axi_master_wstrb,                                     --                                                           .wstrb
			hps_0_h2f_axi_master_wlast                                       => hps_0_h2f_axi_master_wlast,                                     --                                                           .wlast
			hps_0_h2f_axi_master_wvalid                                      => hps_0_h2f_axi_master_wvalid,                                    --                                                           .wvalid
			hps_0_h2f_axi_master_wready                                      => hps_0_h2f_axi_master_wready,                                    --                                                           .wready
			hps_0_h2f_axi_master_bid                                         => hps_0_h2f_axi_master_bid,                                       --                                                           .bid
			hps_0_h2f_axi_master_bresp                                       => hps_0_h2f_axi_master_bresp,                                     --                                                           .bresp
			hps_0_h2f_axi_master_bvalid                                      => hps_0_h2f_axi_master_bvalid,                                    --                                                           .bvalid
			hps_0_h2f_axi_master_bready                                      => hps_0_h2f_axi_master_bready,                                    --                                                           .bready
			hps_0_h2f_axi_master_arid                                        => hps_0_h2f_axi_master_arid,                                      --                                                           .arid
			hps_0_h2f_axi_master_araddr                                      => hps_0_h2f_axi_master_araddr,                                    --                                                           .araddr
			hps_0_h2f_axi_master_arlen                                       => hps_0_h2f_axi_master_arlen,                                     --                                                           .arlen
			hps_0_h2f_axi_master_arsize                                      => hps_0_h2f_axi_master_arsize,                                    --                                                           .arsize
			hps_0_h2f_axi_master_arburst                                     => hps_0_h2f_axi_master_arburst,                                   --                                                           .arburst
			hps_0_h2f_axi_master_arlock                                      => hps_0_h2f_axi_master_arlock,                                    --                                                           .arlock
			hps_0_h2f_axi_master_arcache                                     => hps_0_h2f_axi_master_arcache,                                   --                                                           .arcache
			hps_0_h2f_axi_master_arprot                                      => hps_0_h2f_axi_master_arprot,                                    --                                                           .arprot
			hps_0_h2f_axi_master_arvalid                                     => hps_0_h2f_axi_master_arvalid,                                   --                                                           .arvalid
			hps_0_h2f_axi_master_arready                                     => hps_0_h2f_axi_master_arready,                                   --                                                           .arready
			hps_0_h2f_axi_master_rid                                         => hps_0_h2f_axi_master_rid,                                       --                                                           .rid
			hps_0_h2f_axi_master_rdata                                       => hps_0_h2f_axi_master_rdata,                                     --                                                           .rdata
			hps_0_h2f_axi_master_rresp                                       => hps_0_h2f_axi_master_rresp,                                     --                                                           .rresp
			hps_0_h2f_axi_master_rlast                                       => hps_0_h2f_axi_master_rlast,                                     --                                                           .rlast
			hps_0_h2f_axi_master_rvalid                                      => hps_0_h2f_axi_master_rvalid,                                    --                                                           .rvalid
			hps_0_h2f_axi_master_rready                                      => hps_0_h2f_axi_master_rready,                                    --                                                           .rready
			clk_i_clk_clk                                                    => pll_0_outclk0_clk,                                              --                                                  clk_i_clk.clk
			hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset => rst_controller_002_reset_out_reset,                             -- hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
			sld_hub_controller_system_0_reset_reset_bridge_in_reset_reset    => rst_controller_reset_out_reset,                                 --    sld_hub_controller_system_0_reset_reset_bridge_in_reset.reset
			onchip_memory_nios_arm_s2_address                                => mm_interconnect_1_onchip_memory_nios_arm_s2_address,            --                                  onchip_memory_nios_arm_s2.address
			onchip_memory_nios_arm_s2_write                                  => mm_interconnect_1_onchip_memory_nios_arm_s2_write,              --                                                           .write
			onchip_memory_nios_arm_s2_readdata                               => mm_interconnect_1_onchip_memory_nios_arm_s2_readdata,           --                                                           .readdata
			onchip_memory_nios_arm_s2_writedata                              => mm_interconnect_1_onchip_memory_nios_arm_s2_writedata,          --                                                           .writedata
			onchip_memory_nios_arm_s2_byteenable                             => mm_interconnect_1_onchip_memory_nios_arm_s2_byteenable,         --                                                           .byteenable
			onchip_memory_nios_arm_s2_chipselect                             => mm_interconnect_1_onchip_memory_nios_arm_s2_chipselect,         --                                                           .chipselect
			onchip_memory_nios_arm_s2_clken                                  => mm_interconnect_1_onchip_memory_nios_arm_s2_clken,              --                                                           .clken
			onchip_memory_nios_cpu_s2_address                                => mm_interconnect_1_onchip_memory_nios_cpu_s2_address,            --                                  onchip_memory_nios_cpu_s2.address
			onchip_memory_nios_cpu_s2_write                                  => mm_interconnect_1_onchip_memory_nios_cpu_s2_write,              --                                                           .write
			onchip_memory_nios_cpu_s2_readdata                               => mm_interconnect_1_onchip_memory_nios_cpu_s2_readdata,           --                                                           .readdata
			onchip_memory_nios_cpu_s2_writedata                              => mm_interconnect_1_onchip_memory_nios_cpu_s2_writedata,          --                                                           .writedata
			onchip_memory_nios_cpu_s2_byteenable                             => mm_interconnect_1_onchip_memory_nios_cpu_s2_byteenable,         --                                                           .byteenable
			onchip_memory_nios_cpu_s2_chipselect                             => mm_interconnect_1_onchip_memory_nios_cpu_s2_chipselect,         --                                                           .chipselect
			onchip_memory_nios_cpu_s2_clken                                  => mm_interconnect_1_onchip_memory_nios_cpu_s2_clken,              --                                                           .clken
			sld_hub_controller_system_0_s0_address                           => mm_interconnect_1_sld_hub_controller_system_0_s0_address,       --                             sld_hub_controller_system_0_s0.address
			sld_hub_controller_system_0_s0_write                             => mm_interconnect_1_sld_hub_controller_system_0_s0_write,         --                                                           .write
			sld_hub_controller_system_0_s0_read                              => mm_interconnect_1_sld_hub_controller_system_0_s0_read,          --                                                           .read
			sld_hub_controller_system_0_s0_readdata                          => mm_interconnect_1_sld_hub_controller_system_0_s0_readdata,      --                                                           .readdata
			sld_hub_controller_system_0_s0_writedata                         => mm_interconnect_1_sld_hub_controller_system_0_s0_writedata,     --                                                           .writedata
			sld_hub_controller_system_0_s0_burstcount                        => mm_interconnect_1_sld_hub_controller_system_0_s0_burstcount,    --                                                           .burstcount
			sld_hub_controller_system_0_s0_byteenable                        => mm_interconnect_1_sld_hub_controller_system_0_s0_byteenable,    --                                                           .byteenable
			sld_hub_controller_system_0_s0_readdatavalid                     => mm_interconnect_1_sld_hub_controller_system_0_s0_readdatavalid, --                                                           .readdatavalid
			sld_hub_controller_system_0_s0_waitrequest                       => mm_interconnect_1_sld_hub_controller_system_0_s0_waitrequest,   --                                                           .waitrequest
			sld_hub_controller_system_0_s0_debugaccess                       => mm_interconnect_1_sld_hub_controller_system_0_s0_debugaccess    --                                                           .debugaccess
		);

	irq_mapper : component fluid_board_soc_irq_mapper
		port map (
			clk           => open,                     --       clk.clk
			reset         => open,                     -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq, -- receiver0.irq
			sender_irq    => hps_0_f2h_irq0_irq        --    sender.irq
		);

	irq_mapper_001 : component fluid_board_soc_irq_mapper_001
		port map (
			clk        => open,               --       clk.clk
			reset      => open,               -- clk_reset.reset
			sender_irq => hps_0_f2h_irq1_irq  --    sender.irq
		);

	irq_mapper_002 : component fluid_board_soc_irq_mapper_002
		port map (
			clk            => pll_0_outclk0_clk,                  --        clk.clk
			reset          => rst_controller_001_reset_out_reset, --  clk_reset.reset
			receiver0_irq  => irq_mapper_002_receiver0_irq,       --  receiver0.irq
			receiver1_irq  => irq_mapper_002_receiver1_irq,       --  receiver1.irq
			receiver2_irq  => irq_mapper_002_receiver2_irq,       --  receiver2.irq
			receiver3_irq  => irq_mapper_002_receiver3_irq,       --  receiver3.irq
			receiver4_irq  => irq_mapper_002_receiver4_irq,       --  receiver4.irq
			receiver5_irq  => irq_mapper_002_receiver5_irq,       --  receiver5.irq
			receiver6_irq  => irq_mapper_002_receiver6_irq,       --  receiver6.irq
			receiver7_irq  => irq_mapper_receiver0_irq,           --  receiver7.irq
			receiver8_irq  => irq_mapper_002_receiver8_irq,       --  receiver8.irq
			receiver9_irq  => irq_mapper_002_receiver9_irq,       --  receiver9.irq
			receiver10_irq => irq_mapper_002_receiver10_irq,      -- receiver10.irq
			sender_irq     => nios2_qsys_0_d_irq_irq              --     sender.irq
		);

	rst_controller : component fluid_board_soc_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => hps_0_h2f_reset_reset_ports_inv,    -- reset_in0.reset
			reset_in1      => qsys_reset_reset_n_ports_inv,       -- reset_in1.reset
			clk            => pll_0_outclk0_clk,                  --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_001 : component fluid_board_soc_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => qsys_reset_reset_n_ports_inv,           -- reset_in0.reset
			clk            => pll_0_outclk0_clk,                      --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_001_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_in1      => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_002 : component fluid_board_soc_rst_controller_002
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => hps_0_h2f_reset_reset_ports_inv,    -- reset_in0.reset
			clk            => pll_0_outclk0_clk,                  --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	qsys_reset_reset_n_ports_inv <= not qsys_reset_reset_n;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_pio_reset_nios_s1_write_ports_inv <= not mm_interconnect_0_pio_reset_nios_s1_write;

	mm_interconnect_0_timer_0_s1_write_ports_inv <= not mm_interconnect_0_timer_0_s1_write;

	mm_interconnect_0_timer_1_s1_write_ports_inv <= not mm_interconnect_0_timer_1_s1_write;

	mm_interconnect_0_i2c_master_is1_avalon_slave_0_inv <= not i2c_master_is1_avalon_slave_0_waitrequest;

	mm_interconnect_0_i2c_master_is2_avalon_slave_0_inv <= not i2c_master_is2_avalon_slave_0_waitrequest;

	mm_interconnect_0_i2c_master_is3_avalon_slave_0_inv <= not i2c_master_is3_avalon_slave_0_waitrequest;

	mm_interconnect_0_i2c_master_is4_avalon_slave_0_inv <= not i2c_master_is4_avalon_slave_0_waitrequest;

	mm_interconnect_0_pio_input_s1_write_ports_inv <= not mm_interconnect_0_pio_input_s1_write;

	mm_interconnect_0_pio_output_s1_write_ports_inv <= not mm_interconnect_0_pio_output_s1_write;

	mm_interconnect_0_i2c_master_d_avalon_slave_0_inv <= not i2c_master_d_avalon_slave_0_waitrequest;

	mm_interconnect_0_i2c_master_f_avalon_slave_0_inv <= not i2c_master_f_avalon_slave_0_waitrequest;

	mm_interconnect_0_i2c_master_p_avalon_slave_0_inv <= not i2c_master_p_avalon_slave_0_waitrequest;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	hps_0_h2f_reset_reset_ports_inv <= not hps_0_h2f_reset_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

	pll_0_sys_reset_reset_n <= qsys_reset_reset_n;

	pll_0_sys_clk_clk <= pll_0_outclk0_clk;

end architecture rtl; -- of fluid_board_soc
